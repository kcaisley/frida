* Sampling switch implementation with PMOS/NMOS pair
* Drains and sources connected, gates driven by opposite polarity

*.SCALE METER

.subckt sampswitch vin vout clk clk_b vdd_a vss_a
*.PININFO vin:I vout:O clk:I clk_b:I vdd_a:B vss_a:B

Mp1 vout clk_b vin vdd_a pch_lvt l=60n w=5u m=1
Mn1 vout clk vin vss_a nch_lvt l=60n w=4u m=1

.ends sampswitch
