// Verilog HDL for "basic", "cds_thrualias" "functional"

module cds_thrualias (.thru2(a), .thru1(a));
    inout a;

endmodule
