* ADC Top-level Module - Complete mixed-signal ADC with connectivity between digital and analog blocks

*.BUSDELIMITER [

.SUBCKT adc seq_init seq_samp seq_comp seq_update comp_out en_init en_samp_p en_samp_n en_comp en_update dac_mode dac_diffcaps dac_astate_p[15] dac_astate_p[14] dac_astate_p[13] dac_astate_p[12] dac_astate_p[11] dac_astate_p[10] dac_astate_p[9] dac_astate_p[8] dac_astate_p[7] dac_astate_p[6] dac_astate_p[5] dac_astate_p[4] dac_astate_p[3] dac_astate_p[2] dac_astate_p[1] dac_astate_p[0] dac_bstate_p[15] dac_bstate_p[14] dac_bstate_p[13] dac_bstate_p[12] dac_bstate_p[11] dac_bstate_p[10] dac_bstate_p[9] dac_bstate_p[8] dac_bstate_p[7] dac_bstate_p[6] dac_bstate_p[5] dac_bstate_p[4] dac_bstate_p[3] dac_bstate_p[2] dac_bstate_p[1] dac_bstate_p[0] dac_astate_n[15] dac_astate_n[14] dac_astate_n[13] dac_astate_n[12] dac_astate_n[11] dac_astate_n[10] dac_astate_n[9] dac_astate_n[8] dac_astate_n[7] dac_astate_n[6] dac_astate_n[5] dac_astate_n[4] dac_astate_n[3] dac_astate_n[2] dac_astate_n[1] dac_astate_n[0] dac_bstate_n[15] dac_bstate_n[14] dac_bstate_n[13] dac_bstate_n[12] dac_bstate_n[11] dac_bstate_n[10] dac_bstate_n[9] dac_bstate_n[8] dac_bstate_n[7] dac_bstate_n[6] dac_bstate_n[5] dac_bstate_n[4] dac_bstate_n[3] dac_bstate_n[2] dac_bstate_n[1] dac_bstate_n[0] vin_p vin_n vdd_a vss_a vdd_d vss_d vdd_dac vss_dac
*.PININFO seq_init:I seq_samp:I seq_comp:I seq_update:I comp_out:O en_init:I en_samp_p:I en_samp_n:I en_comp:I en_update:I dac_mode:I dac_diffcaps:I dac_astate_p[15]:I dac_astate_p[14]:I dac_astate_p[13]:I dac_astate_p[12]:I dac_astate_p[11]:I dac_astate_p[10]:I dac_astate_p[9]:I dac_astate_p[8]:I dac_astate_p[7]:I dac_astate_p[6]:I dac_astate_p[5]:I dac_astate_p[4]:I dac_astate_p[3]:I dac_astate_p[2]:I dac_astate_p[1]:I dac_astate_p[0]:I dac_bstate_p[15]:I dac_bstate_p[14]:I dac_bstate_p[13]:I dac_bstate_p[12]:I dac_bstate_p[11]:I dac_bstate_p[10]:I dac_bstate_p[9]:I dac_bstate_p[8]:I dac_bstate_p[7]:I dac_bstate_p[6]:I dac_bstate_p[5]:I dac_bstate_p[4]:I dac_bstate_p[3]:I dac_bstate_p[2]:I dac_bstate_p[1]:I dac_bstate_p[0]:I dac_astate_n[15]:I dac_astate_n[14]:I dac_astate_n[13]:I dac_astate_n[12]:I dac_astate_n[11]:I dac_astate_n[10]:I dac_astate_n[9]:I dac_astate_n[8]:I dac_astate_n[7]:I dac_astate_n[6]:I dac_astate_n[5]:I dac_astate_n[4]:I dac_astate_n[3]:I dac_astate_n[2]:I dac_astate_n[1]:I dac_astate_n[0]:I dac_bstate_n[15]:I dac_bstate_n[14]:I dac_bstate_n[13]:I dac_bstate_n[12]:I dac_bstate_n[11]:I dac_bstate_n[10]:I dac_bstate_n[9]:I dac_bstate_n[8]:I dac_bstate_n[7]:I dac_bstate_n[6]:I dac_bstate_n[5]:I dac_bstate_n[4]:I dac_bstate_n[3]:I dac_bstate_n[2]:I dac_bstate_n[1]:I dac_bstate_n[0]:I vin_p:B vin_n:B vdd_a:B vss_a:B vdd_d:B vss_d:B vdd_dac:B vss_dac:B

* Internal wire declarations
* Digital clock signals
* clk_samp_p clk_samp_p_b clk_samp_n clk_samp_n_b clk_comp
* DAC state signals from digital block (64 bits total)
* dac_state_p_main[15:0] dac_state_p_diff[15:0] dac_state_n_main[15:0] dac_state_n_diff[15:0]
* DAC invert signals from digital block (4 bits total)
* dac_invert_p_main dac_invert_p_diff dac_invert_n_main dac_invert_n_diff
* Capacitor driver outputs (64 bits total)
* dac_drive_botplate_main_p[15:0] dac_drive_botplate_diff_p[15:0]
* dac_drive_botplate_main_n[15:0] dac_drive_botplate_diff_n[15:0]
* Analog voltage signals (vdac_p/vdac_n connect sampswitch, caparray, and comparator)
* vdac_p vdac_n comp_out_p comp_out_n

* Digital block instance
Xadc_digital seq_init seq_samp seq_comp seq_update en_init en_samp_p en_samp_n en_comp en_update dac_mode dac_diffcaps dac_astate_p[15] dac_astate_p[14] dac_astate_p[13] dac_astate_p[12] dac_astate_p[11] dac_astate_p[10] dac_astate_p[9] dac_astate_p[8] dac_astate_p[7] dac_astate_p[6] dac_astate_p[5] dac_astate_p[4] dac_astate_p[3] dac_astate_p[2] dac_astate_p[1] dac_astate_p[0] dac_bstate_p[15] dac_bstate_p[14] dac_bstate_p[13] dac_bstate_p[12] dac_bstate_p[11] dac_bstate_p[10] dac_bstate_p[9] dac_bstate_p[8] dac_bstate_p[7] dac_bstate_p[6] dac_bstate_p[5] dac_bstate_p[4] dac_bstate_p[3] dac_bstate_p[2] dac_bstate_p[1] dac_bstate_p[0] dac_astate_n[15] dac_astate_n[14] dac_astate_n[13] dac_astate_n[12] dac_astate_n[11] dac_astate_n[10] dac_astate_n[9] dac_astate_n[8] dac_astate_n[7] dac_astate_n[6] dac_astate_n[5] dac_astate_n[4] dac_astate_n[3] dac_astate_n[2] dac_astate_n[1] dac_astate_n[0] dac_bstate_n[15] dac_bstate_n[14] dac_bstate_n[13] dac_bstate_n[12] dac_bstate_n[11] dac_bstate_n[10] dac_bstate_n[9] dac_bstate_n[8] dac_bstate_n[7] dac_bstate_n[6] dac_bstate_n[5] dac_bstate_n[4] dac_bstate_n[3] dac_bstate_n[2] dac_bstate_n[1] dac_bstate_n[0] comp_out_p comp_out_n clk_samp_p clk_samp_p_b clk_samp_n clk_samp_n_b clk_comp dac_state_p_main[15] dac_state_p_main[14] dac_state_p_main[13] dac_state_p_main[12] dac_state_p_main[11] dac_state_p_main[10] dac_state_p_main[9] dac_state_p_main[8] dac_state_p_main[7] dac_state_p_main[6] dac_state_p_main[5] dac_state_p_main[4] dac_state_p_main[3] dac_state_p_main[2] dac_state_p_main[1] dac_state_p_main[0] dac_state_p_diff[15] dac_state_p_diff[14] dac_state_p_diff[13] dac_state_p_diff[12] dac_state_p_diff[11] dac_state_p_diff[10] dac_state_p_diff[9] dac_state_p_diff[8] dac_state_p_diff[7] dac_state_p_diff[6] dac_state_p_diff[5] dac_state_p_diff[4] dac_state_p_diff[3] dac_state_p_diff[2] dac_state_p_diff[1] dac_state_p_diff[0] dac_state_n_main[15] dac_state_n_main[14] dac_state_n_main[13] dac_state_n_main[12] dac_state_n_main[11] dac_state_n_main[10] dac_state_n_main[9] dac_state_n_main[8] dac_state_n_main[7] dac_state_n_main[6] dac_state_n_main[5] dac_state_n_main[4] dac_state_n_main[3] dac_state_n_main[2] dac_state_n_main[1] dac_state_n_main[0] dac_state_n_diff[15] dac_state_n_diff[14] dac_state_n_diff[13] dac_state_n_diff[12] dac_state_n_diff[11] dac_state_n_diff[10] dac_state_n_diff[9] dac_state_n_diff[8] dac_state_n_diff[7] dac_state_n_diff[6] dac_state_n_diff[5] dac_state_n_diff[4] dac_state_n_diff[3] dac_state_n_diff[2] dac_state_n_diff[1] dac_state_n_diff[0] dac_invert_p_main dac_invert_p_diff dac_invert_n_main dac_invert_n_diff comp_out vdd_d vss_d / adc_digital

* Four capacitor driver instances
Xcapdriver_p_main dac_state_p_main[15] dac_state_p_main[14] dac_state_p_main[13] dac_state_p_main[12] dac_state_p_main[11] dac_state_p_main[10] dac_state_p_main[9] dac_state_p_main[8] dac_state_p_main[7] dac_state_p_main[6] dac_state_p_main[5] dac_state_p_main[4] dac_state_p_main[3] dac_state_p_main[2] dac_state_p_main[1] dac_state_p_main[0] dac_invert_p_main dac_drive_botplate_main_p[15] dac_drive_botplate_main_p[14] dac_drive_botplate_main_p[13] dac_drive_botplate_main_p[12] dac_drive_botplate_main_p[11] dac_drive_botplate_main_p[10] dac_drive_botplate_main_p[9] dac_drive_botplate_main_p[8] dac_drive_botplate_main_p[7] dac_drive_botplate_main_p[6] dac_drive_botplate_main_p[5] dac_drive_botplate_main_p[4] dac_drive_botplate_main_p[3] dac_drive_botplate_main_p[2] dac_drive_botplate_main_p[1] dac_drive_botplate_main_p[0] vdd_dac vss_dac / capdriver

Xcapdriver_p_diff dac_state_p_diff[15] dac_state_p_diff[14] dac_state_p_diff[13] dac_state_p_diff[12] dac_state_p_diff[11] dac_state_p_diff[10] dac_state_p_diff[9] dac_state_p_diff[8] dac_state_p_diff[7] dac_state_p_diff[6] dac_state_p_diff[5] dac_state_p_diff[4] dac_state_p_diff[3] dac_state_p_diff[2] dac_state_p_diff[1] dac_state_p_diff[0] dac_invert_p_diff dac_drive_botplate_diff_p[15] dac_drive_botplate_diff_p[14] dac_drive_botplate_diff_p[13] dac_drive_botplate_diff_p[12] dac_drive_botplate_diff_p[11] dac_drive_botplate_diff_p[10] dac_drive_botplate_diff_p[9] dac_drive_botplate_diff_p[8] dac_drive_botplate_diff_p[7] dac_drive_botplate_diff_p[6] dac_drive_botplate_diff_p[5] dac_drive_botplate_diff_p[4] dac_drive_botplate_diff_p[3] dac_drive_botplate_diff_p[2] dac_drive_botplate_diff_p[1] dac_drive_botplate_diff_p[0] vdd_dac vss_dac / capdriver

Xcapdriver_n_main dac_state_n_main[15] dac_state_n_main[14] dac_state_n_main[13] dac_state_n_main[12] dac_state_n_main[11] dac_state_n_main[10] dac_state_n_main[9] dac_state_n_main[8] dac_state_n_main[7] dac_state_n_main[6] dac_state_n_main[5] dac_state_n_main[4] dac_state_n_main[3] dac_state_n_main[2] dac_state_n_main[1] dac_state_n_main[0] dac_invert_n_main dac_drive_botplate_main_n[15] dac_drive_botplate_main_n[14] dac_drive_botplate_main_n[13] dac_drive_botplate_main_n[12] dac_drive_botplate_main_n[11] dac_drive_botplate_main_n[10] dac_drive_botplate_main_n[9] dac_drive_botplate_main_n[8] dac_drive_botplate_main_n[7] dac_drive_botplate_main_n[6] dac_drive_botplate_main_n[5] dac_drive_botplate_main_n[4] dac_drive_botplate_main_n[3] dac_drive_botplate_main_n[2] dac_drive_botplate_main_n[1] dac_drive_botplate_main_n[0] vdd_dac vss_dac / capdriver

Xcapdriver_n_diff dac_state_n_diff[15] dac_state_n_diff[14] dac_state_n_diff[13] dac_state_n_diff[12] dac_state_n_diff[11] dac_state_n_diff[10] dac_state_n_diff[9] dac_state_n_diff[8] dac_state_n_diff[7] dac_state_n_diff[6] dac_state_n_diff[5] dac_state_n_diff[4] dac_state_n_diff[3] dac_state_n_diff[2] dac_state_n_diff[1] dac_state_n_diff[0] dac_invert_n_diff dac_drive_botplate_diff_n[15] dac_drive_botplate_diff_n[14] dac_drive_botplate_diff_n[13] dac_drive_botplate_diff_n[12] dac_drive_botplate_diff_n[11] dac_drive_botplate_diff_n[10] dac_drive_botplate_diff_n[9] dac_drive_botplate_diff_n[8] dac_drive_botplate_diff_n[7] dac_drive_botplate_diff_n[6] dac_drive_botplate_diff_n[5] dac_drive_botplate_diff_n[4] dac_drive_botplate_diff_n[3] dac_drive_botplate_diff_n[2] dac_drive_botplate_diff_n[1] dac_drive_botplate_diff_n[0] vdd_dac vss_dac / capdriver

* Two capacitor array instances (cap_shieldplate connected to vss_a)
Xcaparray_p vdac_p vss_a dac_drive_botplate_main_p[15] dac_drive_botplate_main_p[14] dac_drive_botplate_main_p[13] dac_drive_botplate_main_p[12] dac_drive_botplate_main_p[11] dac_drive_botplate_main_p[10] dac_drive_botplate_main_p[9] dac_drive_botplate_main_p[8] dac_drive_botplate_main_p[7] dac_drive_botplate_main_p[6] dac_drive_botplate_main_p[5] dac_drive_botplate_main_p[4] dac_drive_botplate_main_p[3] dac_drive_botplate_main_p[2] dac_drive_botplate_main_p[1] dac_drive_botplate_main_p[0] dac_drive_botplate_diff_p[15] dac_drive_botplate_diff_p[14] dac_drive_botplate_diff_p[13] dac_drive_botplate_diff_p[12] dac_drive_botplate_diff_p[11] dac_drive_botplate_diff_p[10] dac_drive_botplate_diff_p[9] dac_drive_botplate_diff_p[8] dac_drive_botplate_diff_p[7] dac_drive_botplate_diff_p[6] dac_drive_botplate_diff_p[5] dac_drive_botplate_diff_p[4] dac_drive_botplate_diff_p[3] dac_drive_botplate_diff_p[2] dac_drive_botplate_diff_p[1] dac_drive_botplate_diff_p[0] / caparray

Xcaparray_n vdac_n vss_a dac_drive_botplate_main_n[15] dac_drive_botplate_main_n[14] dac_drive_botplate_main_n[13] dac_drive_botplate_main_n[12] dac_drive_botplate_main_n[11] dac_drive_botplate_main_n[10] dac_drive_botplate_main_n[9] dac_drive_botplate_main_n[8] dac_drive_botplate_main_n[7] dac_drive_botplate_main_n[6] dac_drive_botplate_main_n[5] dac_drive_botplate_main_n[4] dac_drive_botplate_main_n[3] dac_drive_botplate_main_n[2] dac_drive_botplate_main_n[1] dac_drive_botplate_main_n[0] dac_drive_botplate_diff_n[15] dac_drive_botplate_diff_n[14] dac_drive_botplate_diff_n[13] dac_drive_botplate_diff_n[12] dac_drive_botplate_diff_n[11] dac_drive_botplate_diff_n[10] dac_drive_botplate_diff_n[9] dac_drive_botplate_diff_n[8] dac_drive_botplate_diff_n[7] dac_drive_botplate_diff_n[6] dac_drive_botplate_diff_n[5] dac_drive_botplate_diff_n[4] dac_drive_botplate_diff_n[3] dac_drive_botplate_diff_n[2] dac_drive_botplate_diff_n[1] dac_drive_botplate_diff_n[0] / caparray

* Two sampling switch instances
Xsampswitch_p vin_p vdac_p clk_samp_p clk_samp_p_b vdd_a vss_a / sampswitch

Xsampswitch_n vin_n vdac_n clk_samp_n clk_samp_n_b vdd_a vss_a / sampswitch

* One comparator instance
Xcomp vdac_p vdac_n comp_out_p comp_out_n clk_comp vdd_a vss_a / comp

.ENDS adc
