VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO c
  CLASS COVER ;
  ORIGIN 0 0 ;
  SIZE 19 BY 19 ;
END c

END LIBRARY