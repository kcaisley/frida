************************************************************************
* auCdl Netlist:
* 
* Library Name:  frida
* Top Cell Name: frida_top
* View Name:     schematic
* Netlisted on:  Oct 16 20:08:09 2025
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: IOlib
* Cell Name:    INVD1_dnw_2_2
* View Name:    schematic
************************************************************************

.SUBCKT INVD1_dnw_2_2 I VDD VSS ZN
*.PININFO I:I ZN:O VDD:B VSS:B
MM0 ZN I VDD VDD pch l=120.0n w=1.04u m=1
MM1 ZN I VSS VSS nch_dnw l=120.0n w=780.0n m=1
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    OPAMP_CMFB_V4_dnw
* View Name:    schematic
************************************************************************

.SUBCKT OPAMP_CMFB_V4_dnw AGND AVDD INN INP OFF OUT VBIAS_OTA
*.PININFO INN:I INP:I OFF:I VBIAS_OTA:I OUT:O AGND:B AVDD:B
MM10 OUT net62 AGND AGND nch_dnw l=1u w=20u m=1
MM16 net14 AGND AGND AGND nch_dnw l=130.0n w=20u m=1
MM9 net14 net56 AGND AGND nch_dnw l=1u w=20u m=1
MM5 net62 net62 AGND AGND nch_dnw l=1u w=20u m=4
MM8 net56 net56 AGND AGND nch_dnw l=1u w=20u m=4
MM17 OUT AGND AGND AGND nch_dnw l=130.0n w=20u m=1
MM15 AVDD AVDD AVDD AVDD pch l=130.0n w=25.0u m=2
MM7 VBIAS_OTA VBIAS_OTA AVDD AVDD pch l=1u w=25.0u m=4
MM0 net20 VBIAS_OTA AVDD AVDD pch l=1u w=25.0u m=8
MM18 VBIAS_OTA VBIAS_OTA VBIAS_OTA AVDD pch l=130.0n w=25.0u m=2
MM3 net62 INP net20 AVDD pch l=1u w=20u m=4
MM12 OUT net14 AVDD AVDD pch l=1u w=20u m=2
MM6 net20 net20 net20 AVDD pch l=130.0n w=20u m=1
MM4 net20 net20 net20 AVDD pch l=130.0n w=20u m=1
MM1 AVDD AVDD AVDD AVDD pch l=130.0n w=20u m=2
MM13 AGND OFF net40 AVDD pch l=130.0n w=2u m=1
MM14 net40 net40 VBIAS_OTA AVDD pch l=1u w=25.0u m=2
MM11 net14 net14 AVDD AVDD pch l=1u w=20u m=2
MM2 net56 INN net20 AVDD pch l=1u w=20u m=4
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    TOP_TX_DUT_v6
* View Name:    schematic
************************************************************************

.SUBCKT TOP_TX_DUT_v6 AGND AVDD AVSS B[0] B[1] B[2] CMFB_IN_N CMFB_IN_P IN 
+ I_DRIVER_EXT OFF OUTN OUTP VBIAS_OTA VREF_CM
*.PININFO B[0]:I B[1]:I B[2]:I CMFB_IN_N:I CMFB_IN_P:I IN:I I_DRIVER_EXT:I 
*.PININFO OFF:I VBIAS_OTA:I VREF_CM:I OUTN:O OUTP:O AGND:B AVDD:B AVSS:B
XR13 net065 net065 rnpolywo l=35.0u w=1u m=1
XR11 net024 net024 rnpolywo l=35.0u w=1u m=1
XR12 net053 net053 rnpolywo l=16.0u w=1u m=1
XR10 net059 net059 rnpolywo l=16.0u w=1u m=1
XR4 net75 I_DRIVER_EXT rnpolywo l=192.000000u w=1u m=1
XR5 net77 I_DRIVER_EXT rnpolywo l=192.000000u w=1u m=1
XR2 net79 I_DRIVER_EXT rnpolywo l=64.0u w=1u m=1
XR20 net84 net83 rnpolywo l=35.0u w=1u m=1
XR19 net83 net82 rnpolywo l=35.0u w=1u m=1
XR18 net82 VREF_CM rnpolywo l=35.0u w=1u m=1
XR16 VREF_CM net80 rnpolywo l=35.0u w=1u m=1
XR15 net80 net067 rnpolywo l=35.0u w=1u m=1
XR14 net067 AGND rnpolywo l=35.0u w=1u m=1
MM24 net0179 AVDD net0190 AGND nch_dnw l=120.0n w=2u m=1
MM2 I_DRIVER_EXT OFF AGND AGND nch_dnw l=130.0n w=2u m=1
MM25 net28 net06 net28 AGND nch_dnw l=4.45u w=4.45u m=6
XI17 B[0] AVDD AGND net74 / INVD1_dnw_2_2
XI16 B[1] AVDD AGND net76 / INVD1_dnw_2_2
XI13 B[2] AVDD AGND net78 / INVD1_dnw_2_2
MM29 net0190 AGND net0179 AVDD pch l=120.0n w=1.2u m=1
MM7 net75 net74 AVDD AVDD pch l=130.0n w=15.0u m=1
MM1 net77 net76 AVDD AVDD pch l=130.0n w=15.0u m=1
MM0 net79 net78 AVDD AVDD pch l=130.0n w=7.5u m=2
MM12 AVDD AVDD AVDD AVDD pch l=200n w=25.0u m=2
MM6 net28 net06 AVDD AVDD pch l=200n w=25.0u m=32
MM10 net84 OFF AVDD AVDD pch l=130.0n w=15.0u m=1
XR8 AGND AGND rppolywo l=1u w=10u m=1
XR7 AGND AGND rppolywo l=1u w=10u m=1
XR6 net40 CMFB_IN_P rppolywo l=15.0u w=10u m=1
XR3 net40 CMFB_IN_N rppolywo l=15.0u w=10u m=1
MM48 AGND AGND OUTN AGND nch_lvt_dnw l=120.0n w=23.0u m=2
MM49 AGND AGND net28 AGND nch_lvt_dnw l=120.0n w=23.0u m=2
MM4 OUTP INN net63 AGND nch_lvt_dnw l=120.0n w=23.0u m=16
MM9 net28 INP OUTP AGND nch_lvt_dnw l=120.0n w=23.0u m=16
MM13 AGND AGND net28 AGND nch_lvt_dnw l=120.0n w=23.0u m=2
MM5 AGND AGND OUTP AGND nch_lvt_dnw l=120.0n w=23.0u m=2
MM3 OUTN INP net63 AGND nch_lvt_dnw l=120.0n w=23.0u m=16
MM8 net28 INN OUTN AGND nch_lvt_dnw l=120.0n w=23.0u m=16
MM15 net63 I_DRIVER_EXT AGND AGND nch_lvt_dnw l=1u w=25.0u m=80
MM14 net63 AGND AGND AGND nch_lvt_dnw l=1u w=25.0u m=8
MM11 I_DRIVER_EXT I_DRIVER_EXT AGND AGND nch_lvt_dnw l=1u w=25.0u m=4
MM16 I_DRIVER_EXT AGND AGND AGND nch_lvt_dnw l=1u w=25.0u m=2
XI21 AGND AVDD VREF_CM net40 OFF net06 VBIAS_OTA / OPAMP_CMFB_V4_dnw
MM46 net0169 IN net0260 AVDD pch l=120.0n w=4.16u m=2
MM45 net0260 OFF AVDD AVDD pch l=120.0n w=4.16u m=2
MM40 INN net0240 AVDD AVDD pch l=120.0n w=2.4u m=16
MM41 INP net0242 AVDD AVDD pch l=120.0n w=2.4u m=16
MM39 net0242 net0230 AVDD AVDD pch l=120.0n w=2.4u m=8
MM38 net0240 net0228 AVDD AVDD pch l=120.0n w=2.4u m=8
MM33 net0230 net0218 AVDD AVDD pch l=120.0n w=2.4u m=4
MM32 net0228 net0216 AVDD AVDD pch l=120.0n w=2.4u m=4
MM28 net0218 net0206 AVDD AVDD pch l=120.0n w=2.4u m=2
MM27 net0216 net0204 AVDD AVDD pch l=120.0n w=2.4u m=2
MM22 net0204 net0190 AVDD AVDD pch l=120.0n w=2.4u m=1
MM21 net0206 net0192 AVDD AVDD pch l=120.0n w=2.4u m=1
MM19 net0192 net0179 AVDD AVDD pch l=120.0n w=2.4u m=1
MM17 net0179 net0169 AVDD AVDD pch l=120.0n w=2.4u m=4
MM47 net0169 IN AGND AGND nch_dnw l=120.0n w=3.12u m=2
MM44 net0169 OFF AGND AGND nch_dnw l=120.0n w=3.12u m=2
MM43 INP net0242 AGND AGND nch_dnw l=120.0n w=800n m=16
MM42 INN net0240 AGND AGND nch_dnw l=120.0n w=800n m=16
MM37 net0242 net0230 AGND AGND nch_dnw l=120.0n w=800n m=8
MM36 net0240 net0228 AGND AGND nch_dnw l=120.0n w=800n m=8
MM35 net0230 net0218 AGND AGND nch_dnw l=120.0n w=800n m=4
MM34 net0228 net0216 AGND AGND nch_dnw l=120.0n w=800n m=4
MM31 net0218 net0206 AGND AGND nch_dnw l=120.0n w=800n m=2
MM30 net0216 net0204 AGND AGND nch_dnw l=120.0n w=800n m=2
MM26 net0204 net0190 AGND AGND nch_dnw l=120.0n w=800n m=1
MM23 net0206 net0192 AGND AGND nch_dnw l=120.0n w=800n m=1
MM20 net0192 net0179 AGND AGND nch_dnw l=120.0n w=800n m=1
MM18 net0179 net0169 AGND AGND nch_dnw l=120.0n w=800n m=4
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    SF_1V2_CDM
* View Name:    schematic
************************************************************************

.SUBCKT SF_1V2_CDM IO Internal VDD VDDPST VSS VSSPST
*.PININFO IO:B Internal:B VDD:B VDDPST:B VSS:B VSSPST:B
MM0 Internal VSSPST VSSPST VSSPST nch l=6e-08 w=6.06e-05 m=1
MM2 Internal VDDPST VDDPST VDDPST pch l=1e-07 w=5.672e-05 m=1
DD4 N0 VSSPST ndio area=5.45292e-11 pj=4e-05 m=1
DD6 VSSPST IO ndio area=5.20506e-11 pj=4e-05 m=1
DD7 VSSPST VDDPST ndio area=5.45292e-11 pj=4e-05 m=1
DD8 IO N1 pdio area=3.55266e-11 pj=4e-05 m=1
DD10 N1 N2 pdio area=5.20506e-11 pj=4e-05 m=1
DD11 N2 N3 pdio area=2.60253e-11 pj=4e-05 m=1
DD12 N3 VSSPST pdio area=2.60253e-11 pj=4e-05 m=1
DD13 N4 VSSPST pdio area=2.60253e-11 pj=4e-05 m=1
DD14 N5 N4 pdio area=2.60253e-11 pj=4e-05 m=1
DD16 N1 N5 pdio area=5.20506e-11 pj=4e-05 m=1
DD17 N1 VDDPST pdio area=3.55266e-11 pj=4e-05 m=1
DD18 VDDPST N1 pdio area=3.55266e-11 pj=4e-05 m=1
XR19 Internal IO rppolywo l=1.1e-06 w=3.8e-05 m=1
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    PASSIVE_CUP_pad
* View Name:    schematic
************************************************************************

.SUBCKT PASSIVE_CUP_pad I O PAD VDD VDDPST VSS VSSPST
*.PININFO I:I O:O PAD:B VDD:B VDDPST:B VSS:B VSSPST:B
*.CONNECT I PAD 
XI3 PAD O VDD VDDPST VSS VSSPST / SF_1V2_CDM
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    LVDS_TX_CUP_pad
* View Name:    schematic
************************************************************************

.SUBCKT LVDS_TX_CUP_pad DS[2] DS[1] DS[0] EN_B I PAD_N PAD_P VDD VDDPST VSS 
+ VSSPST
*.PININFO DS[2]:I DS[1]:I DS[0]:I EN_B:I I:I PAD_N:O PAD_P:O VDD:B VDDPST:B 
*.PININFO VSS:B VSSPST:B
XI0 VSSPST VDDPST VSS DS[0] DS[1] DS[2] net15 net16 I net14 EN_B PAD_N PAD_P 
+ net11 net10 / TOP_TX_DUT_v6
XI8 net018 net15 PAD_N VDD VDDPST VSS VSSPST / PASSIVE_CUP_pad
XI11 net017 net16 PAD_P VDD VDDPST VSS VSSPST / PASSIVE_CUP_pad
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    TOP_RX_DUT_v2
* View Name:    schematic
************************************************************************

.SUBCKT TOP_RX_DUT_v2 AVDD AVSS INN INP OFF OUT_RX
*.PININFO INN:I INP:I OFF:I OUT_RX:O AVDD:B AVSS:B
MM13 net0105 net0105 AVDD AVDD pch_lvt l=120.0n w=6u m=1
MM19 net069 OUTN_2 AVDD AVDD pch_lvt l=120.0n w=6u m=1
MM29 net075 AVDD AVDD AVDD pch_lvt l=120.0n w=12.5u m=1
MM28 net075 AVDD AVDD AVDD pch_lvt l=120.0n w=12.5u m=1
MM50 SOURCE net077 AVDD AVDD pch_lvt l=200n w=22.0u m=40
MM27 net075 INP SOURCE AVDD pch_lvt l=120.0n w=12.5u m=2
MM16 OUTN_2 OUTP_2 AVDD AVDD pch_lvt l=120.0n w=6u m=1
MM30 net076 INN SOURCE AVDD pch_lvt l=120.0n w=12.5u m=2
MM44 net017 net017 net077 AVDD pch_lvt l=1u w=6.5u m=1
MM18 OUTN_2 OUTN_2 AVDD AVDD pch_lvt l=120.0n w=6u m=1
MM2 AVDD net077 AVDD AVDD pch_lvt l=200n w=22.0u m=1
MM1 AVDD net077 AVDD AVDD pch_lvt l=200n w=22.0u m=1
MM15 OUTP_2 OUTN_2 AVDD AVDD pch_lvt l=120.0n w=6u m=1
MM10 net0125 net0105 AVDD AVDD pch_lvt l=120.0n w=6u m=1
MM49 net077 net077 AVDD AVDD pch_lvt l=200n w=22.0u m=4
MM20 net0125 OUTP_2 AVDD AVDD pch_lvt l=120.0n w=6u m=1
MM17 OUTP_2 OUTP_2 AVDD AVDD pch_lvt l=120.0n w=6u m=1
MM35 net0128 net0125 AVDD AVDD pch l=130.0n w=400n m=2
MM34 net0105 nOFF AVDD AVDD pch l=130.0n w=1u m=1
MMU1-M_u3 nOFF OFF AVDD AVDD pch l=120.0n w=1.04u m=1
MM39 OUT_RX net0128 AVDD AVDD pch l=130.0n w=400n m=4
MM0 net016 OFF AVDD AVDD pch l=130.0n w=1u m=1
MM8 net0105 net076 AVSS AVSS nch_lvt_dnw l=120.0n w=6u m=1
MM9 net0125 net075 AVSS AVSS nch_lvt_dnw l=120.0n w=6u m=1
MM23 net076 net075 AVSS AVSS nch_lvt_dnw l=120.0n w=3u m=1
MM26 net076 net076 AVSS AVSS nch_lvt_dnw l=120.0n w=3u m=1
MM12 OUTP_2 INP I_OUT AVSS nch_lvt_dnw l=120.0n w=10u m=1
MM3 I_OUT net013 AVSS AVSS nch_lvt_dnw l=200n w=22.0u m=40
MM6 net075 net075 AVSS AVSS nch_lvt_dnw l=120.0n w=3u m=1
MM21 net069 net069 AVSS AVSS nch_lvt_dnw l=120.0n w=2u m=1
MM11 net075 net076 AVSS AVSS nch_lvt_dnw l=120.0n w=3u m=1
MM4 AVSS net013 AVSS AVSS nch_lvt_dnw l=200n w=22.0u m=1
MM22 net0125 net069 AVSS AVSS nch_lvt_dnw l=120.0n w=2u m=1
MM5 AVSS net013 AVSS AVSS nch_lvt_dnw l=200n w=22.0u m=1
MM14 OUTN_2 INN I_OUT AVSS nch_lvt_dnw l=120.0n w=10u m=1
MM24 net013 net013 AVSS AVSS nch_lvt_dnw l=200n w=22.0u m=4
MM48 net017 nOFF AVSS AVSS nch_dnw l=130.0n w=1u m=1
MM38 OUT_RX net0128 AVSS AVSS nch_dnw l=130.0n w=200n m=4
MM36 net0128 net0125 AVSS AVSS nch_dnw l=130.0n w=200n m=2
MM33 net069 OFF AVSS AVSS nch_dnw l=130.0n w=1u m=1
MMU1-M_u2 nOFF OFF AVSS AVSS nch_dnw l=120.0n w=780.0n m=1
MM25 net016 net016 net013 AVSS nch_dnw l=1u w=2u m=1
MM7 net0125 OFF AVSS AVSS nch_dnw l=130.0n w=1u m=1
XR15 INP AVDD rppolywo l=75.55u w=3u m=1
XR12 AVDD INN rppolywo l=75.55u w=3u m=1
XR10 INN AVSS rppolywo l=35.26u w=5u m=1
XR16 AVSS INP rppolywo l=32.71u w=5u m=1
.ENDS

************************************************************************
* Library Name: tcbn65lp_dnw
* Cell Name:    DCAP64
* View Name:    schematic
************************************************************************

.SUBCKT DCAP64 VDD VSS
*.PININFO VDD:B VSS:B
MMI54 VDD net11 VDD VDD pch l=915.00n w=430.0n m=1
MM_u1 net67 net11 VDD VDD pch l=60n w=390.0n m=1
MMI56 VDD net11 VDD VDD pch l=915.00n w=430.0n m=1
MMI55 VDD net11 VDD VDD pch l=915.00n w=430.0n m=1
MMI39 VDD net11 VDD VDD pch l=915.00n w=430.0n m=1
MMI57 VDD net11 VDD VDD pch l=915.00n w=430.0n m=1
MMI58 VDD net11 VDD VDD pch l=915.00n w=430.0n m=1
MMI59 VDD net11 VDD VDD pch l=915.00n w=430.0n m=1
MMI53 VDD net11 VDD VDD pch l=915.00n w=430.0n m=1
MMI50 VDD net11 VDD VDD pch l=915.00n w=430.0n m=1
MMI52 VDD net11 VDD VDD pch l=915.00n w=430.0n m=1
MMI51 VDD net11 VDD VDD pch l=915.00n w=430.0n m=1
MMI64 VSS net67 VSS VSS nch_dnw l=915.00n w=300n m=1
MMI65 VSS net67 VSS VSS nch_dnw l=915.00n w=300n m=1
MMI62 VSS net67 VSS VSS nch_dnw l=915.00n w=300n m=1
MMI67 VSS net67 VSS VSS nch_dnw l=915.00n w=300n m=1
MMI68 VSS net67 VSS VSS nch_dnw l=915.00n w=300n m=1
MMI60 VSS net67 VSS VSS nch_dnw l=915.00n w=300n m=1
MMI66 VSS net67 VSS VSS nch_dnw l=915.00n w=300n m=1
MMI69 VSS net67 VSS VSS nch_dnw l=915.00n w=300n m=1
MMI49 VSS net67 VSS VSS nch_dnw l=915.00n w=300n m=1
MMI61 VSS net67 VSS VSS nch_dnw l=915.00n w=300n m=1
MM_u2 net11 net67 VSS VSS nch_dnw l=60n w=300n m=1
MMI63 VSS net67 VSS VSS nch_dnw l=915.00n w=300n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lp_dnw
* Cell Name:    CKBD24
* View Name:    schematic
************************************************************************

.SUBCKT CKBD24 I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
DDI3 VSS I ndio area=6.6e-14 pj=1.18e-06 m=1
MMU21_12 Z net5 VDD VDD pch l=60n w=520.0n m=1
MM_u3_4 net5 I VDD VDD pch l=60n w=520.0n m=1
MMU21_15 Z net5 VDD VDD pch l=60n w=520.0n m=1
MMU21_7 Z net5 VDD VDD pch l=60n w=520.0n m=1
MMU21_0 Z net5 VDD VDD pch l=60n w=520.0n m=1
MMU21_17 Z net5 VDD VDD pch l=60n w=520.0n m=1
MMU21_1 Z net5 VDD VDD pch l=60n w=520.0n m=1
MMU21_11 Z net5 VDD VDD pch l=60n w=520.0n m=1
MMU21_16 Z net5 VDD VDD pch l=60n w=520.0n m=1
MMU21_5 Z net5 VDD VDD pch l=60n w=520.0n m=1
MMU21_19 Z net5 VDD VDD pch l=60n w=520.0n m=1
MM_u3_3 net5 I VDD VDD pch l=60n w=520.0n m=1
MM_u3_5 net5 I VDD VDD pch l=60n w=520.0n m=1
MM_u3_0 net5 I VDD VDD pch l=60n w=520.0n m=1
MMU21_23 Z net5 VDD VDD pch l=60n w=520.0n m=1
MMU21_10 Z net5 VDD VDD pch l=60n w=520.0n m=1
MMU21_13 Z net5 VDD VDD pch l=60n w=520.0n m=1
MMU21_3 Z net5 VDD VDD pch l=60n w=520.0n m=1
MMU21_4 Z net5 VDD VDD pch l=60n w=520.0n m=1
MM_u3_2 net5 I VDD VDD pch l=60n w=520.0n m=1
MMU21_22 Z net5 VDD VDD pch l=60n w=520.0n m=1
MMU21_6 Z net5 VDD VDD pch l=60n w=520.0n m=1
MMU21_21 Z net5 VDD VDD pch l=60n w=520.0n m=1
MMU21_18 Z net5 VDD VDD pch l=60n w=520.0n m=1
MMU21_9 Z net5 VDD VDD pch l=60n w=520.0n m=1
MMU21_20 Z net5 VDD VDD pch l=60n w=520.0n m=1
MMU21_8 Z net5 VDD VDD pch l=60n w=520.0n m=1
MM_u3_1 net5 I VDD VDD pch l=60n w=520.0n m=1
MMU21_2 Z net5 VDD VDD pch l=60n w=520.0n m=1
MM_u3_6 net5 I VDD VDD pch l=60n w=520.0n m=1
MMU21_14 Z net5 VDD VDD pch l=60n w=520.0n m=1
MM_u15 net5 I VSS VSS nch_dnw l=60n w=2.1u m=1
MMU23 Z net5 VSS VSS nch_dnw l=60n w=7.35u m=1
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    LVDS_RX_CUP_pad
* View Name:    schematic
************************************************************************

.SUBCKT LVDS_RX_CUP_pad EN_B O PAD_N PAD_P VDD VDDPST VSS VSSPST
*.PININFO EN_B:I PAD_N:I PAD_P:I O:O VDD:B VDDPST:B VSS:B VSSPST:B
XI0 VDDPST VSSPST net15 net12 EN_B net011 / TOP_RX_DUT_v2
XI5 VDDPST VSSPST / DCAP64
XI1 net011 VDDPST VSSPST O / CKBD24
XI8 net014 net15 PAD_N VDD VDDPST VSS VSSPST / PASSIVE_CUP_pad
XI9 net013 net12 PAD_P VDD VDDPST VSS VSSPST / PASSIVE_CUP_pad
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    DNW_DEL0
* View Name:    schematic
************************************************************************

.SUBCKT DNW_DEL0 I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
MMI2-M_u3 Z net11 VDD VDD pch l=60n w=520.0n m=1
MMU5-M_u3 net25 net5 VDD VDD pch l=600n w=520.0n m=1
MMI1-M_u3 net5 I VDD VDD pch l=60n w=520.0n m=1
MMU7-M_u3 net11 net25 VDD VDD pch l=600n w=520.0n m=1
MM3 Z net11 VSS VSS nch_dnw l=60n w=390.0n m=1
MM2 net5 I VSS VSS nch_dnw l=60n w=390.0n m=1
MM1 net25 net5 VSS VSS nch_dnw l=600n w=390.0n m=1
MM0 net11 net25 VSS VSS nch_dnw l=600n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    DNW_DEL015
* View Name:    schematic
************************************************************************

.SUBCKT DNW_DEL015 I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
MMI2-M_u3 Z net13 VDD VDD pch l=60n w=520.0n m=1
MMI20 net57 net9 VDD VDD pch l=60n w=520.0n m=1
MMI23 net13 net9 net25 VDD pch l=60n w=520.0n m=1
MMI1-M_u3 net5 I VDD VDD pch l=60n w=520.0n m=1
MMI21 net25 net9 net57 VDD pch l=60n w=520.0n m=1
MMI32 net9 net5 net44 VDD pch l=60n w=520.0n m=1
MMI31 net44 net5 net33 VDD pch l=60n w=520.0n m=1
MMI7 net33 net5 VDD VDD pch l=60n w=520.0n m=1
MM7 net44 net5 net17 VSS nch_dnw l=60n w=390.0n m=1
MM6 net5 I VSS VSS nch_dnw l=60n w=390.0n m=1
MM5 net9 net5 net44 VSS nch_dnw l=60n w=390.0n m=1
MM4 net13 net9 net25 VSS nch_dnw l=60n w=390.0n m=1
MM3 net17 net5 VSS VSS nch_dnw l=60n w=390.0n m=1
MM2 net28 net9 VSS VSS nch_dnw l=60n w=390.0n m=1
MM1 net25 net9 net28 VSS nch_dnw l=60n w=390.0n m=1
MM0 Z net13 VSS VSS nch_dnw l=60n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    DNW_INR2D2
* View Name:    schematic
************************************************************************

.SUBCKT DNW_INR2D2 A1 B1 VDD VSS ZN
*.PININFO A1:I B1:I ZN:O VDD:B VSS:B
MMU6-M_u3 net5 A1 VDD VDD pch l=60n w=520.0n m=1
MMU1_0-M_u2 ZN B1 net36 VDD pch l=60n w=520.0n m=1
MMU1_0-M_u1 net36 net5 VDD VDD pch l=60n w=520.0n m=1
MMU1_1-M_u1 net25 net5 VDD VDD pch l=60n w=520.0n m=1
MMU1_1-M_u2 ZN B1 net25 VDD pch l=60n w=520.0n m=1
MM4 ZN B1 VSS VSS nch_dnw l=60n w=390.0n m=1
MM3 net5 A1 VSS VSS nch_dnw l=60n w=390.0n m=1
MM2 ZN net5 VSS VSS nch_dnw l=60n w=390.0n m=1
MM1 ZN net5 VSS VSS nch_dnw l=60n w=390.0n m=1
MM0 ZN B1 VSS VSS nch_dnw l=60n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    DNW_INVD1
* View Name:    schematic
************************************************************************

.SUBCKT DNW_INVD1 I VDD VSS ZN
*.PININFO I:I ZN:O VDD:B VSS:B
MMU1-M_u3 ZN I VDD VDD pch l=60n w=520.0n m=1
MM0 ZN I VSS VSS nch_dnw l=60n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    DNW_BUFFD2
* View Name:    schematic
************************************************************************

.SUBCKT DNW_BUFFD2 I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
MM_u3_0-M_u3 Z net11 VDD VDD pch l=60n w=520.0n m=1
MM_u3_1-M_u3 Z net11 VDD VDD pch l=60n w=520.0n m=1
MM_u2-M_u3 net11 I VDD VDD pch l=60n w=520.0n m=1
MM2 Z net11 VSS VSS nch_dnw l=60n w=390.0n m=1
MM1 net11 I VSS VSS nch_dnw l=60n w=390.0n m=1
MM0 Z net11 VSS VSS nch_dnw l=60n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    DNW_NR2D1
* View Name:    schematic
************************************************************************

.SUBCKT DNW_NR2D1 A1 A2 VDD VSS ZN
*.PININFO A1:I A2:I ZN:O VDD:B VSS:B
MMI1-M_u1 net13 A2 VDD VDD pch l=60n w=520.0n m=1
MMI1-M_u2 ZN A1 net13 VDD pch l=60n w=520.0n m=1
MM1 ZN A1 VSS VSS nch_dnw l=60n w=390.0n m=1
MM0 ZN A2 VSS VSS nch_dnw l=60n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    DNW_ND2D1
* View Name:    schematic
************************************************************************

.SUBCKT DNW_ND2D1 A1 A2 VDD VSS ZN
*.PININFO A1:I A2:I ZN:O VDD:B VSS:B
MMI1-M_u1 ZN A1 VDD VDD pch l=60n w=520.0n m=1
MMI1-M_u2 ZN A2 VDD VDD pch l=60n w=520.0n m=1
MM1 net1 A2 VSS VSS nch_dnw l=60n w=390.0n m=1
MM0 ZN A1 net1 VSS nch_dnw l=60n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    PAD_SchmittTrigger
* View Name:    schematic
************************************************************************

.SUBCKT PAD_SchmittTrigger A DS IO Internal OUT_EN PEN UD VDDPST VSSPST Z Z_h
*.PININFO A:I DS:I OUT_EN:I PEN:I UD:I VDDPST:I VSSPST:I Z:O Z_h:O IO:B 
*.PININFO Internal:B
XI84 net226 VDDPST VSSPST net235 / DNW_DEL0
XI83 net229 VDDPST VSSPST net236 / DNW_DEL0
XI94 net213 VDDPST VSSPST net212 / DNW_DEL015
XI93 net212 VDDPST VSSPST net217 / DNW_DEL015
XI92 net217 VDDPST VSSPST net078 / DNW_DEL015
XI85 net020 VDDPST VSSPST net215 / DNW_DEL015
XI90 net223 VDDPST VSSPST net226 / DNW_DEL015
XI87 net219 VDDPST VSSPST net222 / DNW_DEL015
XI88 net222 VDDPST VSSPST net075 / DNW_DEL015
XI89 net075 VDDPST VSSPST net229 / DNW_DEL015
XI86 net215 VDDPST VSSPST net219 / DNW_DEL015
XI91 net078 VDDPST VSSPST net223 / DNW_DEL015
XI107 PEN UD VDDPST VSSPST net071 / DNW_INR2D2
XI108 net090 VDDPST VSSPST Z_h / DNW_INVD1
XI76 net058 VDDPST VSSPST net230 / DNW_INVD1
XI74 net250 VDDPST VSSPST net213 / DNW_INVD1
XI78 OUT_EN VDDPST VSSPST net251 / DNW_INVD1
XI75 net057 VDDPST VSSPST net227 / DNW_INVD1
XI77 DS VDDPST VSSPST net234 / DNW_INVD1
XI73 net249 VDDPST VSSPST net020 / DNW_INVD1
MM16 VSSPST net090 net066 VDDPST pch l=60n w=1.55u m=1
MM10 net090 Internal net066 VDDPST pch l=60n w=1.55u m=1
MM9 net066 Internal VDDPST VDDPST pch l=60n w=1.55u m=1
MM7 Internal net070 net069 VDDPST pch l=60n w=1.55u m=1
MM34 IO net237 VDDPST VDDPST pch l=60n w=1.55u m=36
MM32 IO net239 VDDPST VDDPST pch l=60n w=1.55u m=36
MM30 IO net241 VDDPST VDDPST pch l=60n w=1.55u m=8
MM20 IO net243 VDDPST VDDPST pch l=60n w=1.55u m=8
MM15 IO net245 VDDPST VDDPST pch l=60n w=1.55u m=6
MM14 IO net247 VDDPST VDDPST pch l=60n w=1.55u m=6
MM13 IO net209 VDDPST VDDPST pch l=60n w=1.55u m=6
XI80 net206 VDDPST VSSPST net250 / DNW_BUFFD2
XI81 net251 VDDPST VSSPST net232 / DNW_BUFFD2
XI79 net209 VDDPST VSSPST net249 / DNW_BUFFD2
XI82 Internal VDDPST VSSPST Z / DNW_BUFFD2
XI97 A net232 VDDPST VSSPST net206 / DNW_NR2D1
XI98 net234 net213 VDDPST VSSPST net057 / DNW_NR2D1
XI103 net213 net217 VDDPST VSSPST net246 / DNW_NR2D1
XI99 net227 net235 VDDPST VSSPST net238 / DNW_NR2D1
XI100 net227 net226 VDDPST VSSPST net240 / DNW_NR2D1
XI101 net213 net223 VDDPST VSSPST net242 / DNW_NR2D1
XI104 net213 net212 VDDPST VSSPST net248 / DNW_NR2D1
XI102 net213 net078 VDDPST VSSPST net244 / DNW_NR2D1
MM17 VDDPST net090 net025 VSSPST nch_dnw l=60n w=700n m=1
MM12 net025 Internal VSSPST VSSPST nch_dnw l=60n w=700n m=1
MM11 net090 Internal net025 VSSPST nch_dnw l=60n w=700n m=1
MM8 Internal net071 net092 VSSPST nch_dnw l=60n w=700n m=1
MM2 IO net246 VSSPST VSSPST nch_dnw l=60n w=700n m=6
MM1 IO net248 VSSPST VSSPST nch_dnw l=60n w=700n m=6
MM0 IO net206 VSSPST VSSPST nch_dnw l=60n w=700n m=6
MM5 IO net240 VSSPST VSSPST nch_dnw l=60n w=700n m=36
MM6 IO net238 VSSPST VSSPST nch_dnw l=60n w=700n m=36
MM3 IO net244 VSSPST VSSPST nch_dnw l=60n w=700n m=8
MM4 IO net242 VSSPST VSSPST nch_dnw l=60n w=700n m=8
DD0 Internal VDDPST pdio area=4.095e-10 pj=8.1e-05 m=1
XR0 VSSPST net092 rppolywo l=55.825u w=1u m=1
XR1 VDDPST net069 rppolywo l=55.825u w=1u m=1
XI106 PEN UD VDDPST VSSPST net070 / DNW_ND2D1
XI65 A OUT_EN VDDPST VSSPST net209 / DNW_ND2D1
XI66 DS net020 VDDPST VSSPST net058 / DNW_ND2D1
XI67 net020 net215 VDDPST VSSPST net247 / DNW_ND2D1
XI68 net020 net222 VDDPST VSSPST net243 / DNW_ND2D1
XI69 net020 net219 VDDPST VSSPST net245 / DNW_ND2D1
XI70 net020 net075 VDDPST VSSPST net241 / DNW_ND2D1
XI71 net230 net229 VDDPST VSSPST net239 / DNW_ND2D1
XI72 net230 net236 VDDPST VSSPST net237 / DNW_ND2D1
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    CMOS_IO_CUP_pad
* View Name:    schematic
************************************************************************

.SUBCKT CMOS_IO_CUP_pad A DS OUT_EN PAD PEN UD_B VDD VDDPST VSS VSSPST Z Z_h
*.PININFO A:I DS:I OUT_EN:I PEN:I UD_B:I Z:O Z_h:O PAD:B VDD:B VDDPST:B VSS:B 
*.PININFO VSSPST:B
XI13 A DS PAD Internal OUT_EN PEN UD_B VDDPST VSSPST Z Z_h / PAD_SchmittTrigger
XI3 PAD Internal VDD VDDPST VSS VSSPST / SF_1V2_CDM
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    SF_1V2_POWER_CLAMP_IO_SUPPLY
* View Name:    schematic
************************************************************************

.SUBCKT SF_1V2_POWER_CLAMP_IO_SUPPLY VDD VDDPST VSS VSSPST
*.PININFO VDD:B VDDPST:B VSS:B VSSPST:B
DD0 N0 VSSPST ndio area=5.45292e-11 pj=4e-05 m=1
DD1 VSSPST VDDPST ndio area=5.45292e-11 pj=4e-05 m=1
DD2 N1 VSSPST pdio area=2.60253e-11 pj=4e-05 m=1
DD3 N2 N1 pdio area=2.60253e-11 pj=4e-05 m=1
DD5 N3 N2 pdio area=5.20506e-11 pj=4e-05 m=1
DD6 VDDPST N3 pdio area=3.55266e-11 pj=4e-05 m=1
DD7 VSSPST VSS pdio area=3.55266e-11 pj=4e-05 m=1
DD8 VSS VSSPST pdio area=3.55266e-11 pj=4e-05 m=1
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    POWER_CUP_pad
* View Name:    schematic
************************************************************************

.SUBCKT POWER_CUP_pad VDD VDDPST VSS VSSPST
*.PININFO VDD:B VDDPST:B VSS:B VSSPST:B
XI0 VDD VDDPST VSS VSSPST / SF_1V2_POWER_CLAMP_IO_SUPPLY
XR0[9] VDD VDDPST rm2 l=2u w=1.2u m=1
XR0[8] VDD VDDPST rm2 l=2u w=1.2u m=1
XR0[7] VDD VDDPST rm2 l=2u w=1.2u m=1
XR0[6] VDD VDDPST rm2 l=2u w=1.2u m=1
XR0[5] VDD VDDPST rm2 l=2u w=1.2u m=1
XR0[4] VDD VDDPST rm2 l=2u w=1.2u m=1
XR0[3] VDD VDDPST rm2 l=2u w=1.2u m=1
XR0[2] VDD VDDPST rm2 l=2u w=1.2u m=1
XR0[1] VDD VDDPST rm2 l=2u w=1.2u m=1
XR0[0] VDD VDDPST rm2 l=2u w=1.2u m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    TIELLVT
* View Name:    schematic
************************************************************************

.SUBCKT TIELLVT VDD VSS ZN
*.PININFO ZN:O VDD:B VSS:B
MM_u2 ZN net5 VSS VSS nch_lvt l=60n w=410.0n m=1
MM_u1 net5 net5 VDD VDD pch_lvt l=60n w=540.0n m=1
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    SF_1V2_POWER_CLAMP_IO_GROUND
* View Name:    schematic
************************************************************************

.SUBCKT SF_1V2_POWER_CLAMP_IO_GROUND VDD VDDPST VSS VSSPST
*.PININFO VDD:B VDDPST:B VSS:B VSSPST:B
DD0 N0 VSSPST ndio area=5.45292e-11 pj=4e-05 m=1
DD1 VSSPST VDDPST ndio area=5.45292e-11 pj=4e-05 m=1
DD2 N1 VSSPST pdio area=2.60253e-11 pj=4e-05 m=1
DD3 N2 N1 pdio area=2.60253e-11 pj=4e-05 m=1
DD5 N3 N2 pdio area=5.20506e-11 pj=4e-05 m=1
DD6 VDDPST N3 pdio area=3.55266e-11 pj=4e-05 m=1
DD7 VSSPST VSS pdio area=3.55266e-11 pj=4e-05 m=1
DD8 VSS VSSPST pdio area=3.55266e-11 pj=4e-05 m=1
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    GROUND_CUP_pad
* View Name:    schematic
************************************************************************

.SUBCKT GROUND_CUP_pad VDD VDDPST VSS VSSPST
*.PININFO VDD:B VDDPST:B VSS:B VSSPST:B
XI0 VDD VDDPST VSS VSSPST / SF_1V2_POWER_CLAMP_IO_GROUND
.ENDS

************************************************************************
* Library Name: tcbn65lp_dnw
* Cell Name:    DCAP32
* View Name:    schematic
************************************************************************

.SUBCKT DCAP32 VDD VSS
*.PININFO VDD:B VSS:B
MMI33 VDD net5 VDD VDD pch l=975.00n w=430.0n m=1
MM_u1 net11 net5 VDD VDD pch l=60n w=390.0n m=1
MMI34 VDD net5 VDD VDD pch l=975.00n w=430.0n m=1
MMI35 VDD net5 VDD VDD pch l=975.00n w=430.0n m=1
MMI32 VDD net5 VDD VDD pch l=975.00n w=430.0n m=1
MMI26 VDD net5 VDD VDD pch l=975.00n w=430.0n m=1
MMI38 VSS net11 VSS VSS nch_dnw l=975.00n w=300n m=1
MMI6 VSS net11 VSS VSS nch_dnw l=975.00n w=300n m=1
MMI39 VSS net11 VSS VSS nch_dnw l=975.00n w=300n m=1
MMI37 VSS net11 VSS VSS nch_dnw l=975.00n w=300n m=1
MM_u2 net5 net11 VSS VSS nch_dnw l=60n w=300n m=1
MMI36 VSS net11 VSS VSS nch_dnw l=975.00n w=300n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lp_dnw
* Cell Name:    DCAP16
* View Name:    schematic
************************************************************************

.SUBCKT DCAP16 VDD VSS
*.PININFO VDD:B VSS:B
MMI3 VDD net5 VDD VDD pch l=690.0n w=430.0n m=1
MMI6 VDD net5 VDD VDD pch l=690.0n w=430.0n m=1
MM_u1 net11 net5 VDD VDD pch l=60n w=390.0n m=1
MMI5 VDD net5 VDD VDD pch l=690.0n w=430.0n m=1
MMI4 VSS net11 VSS VSS nch_dnw l=690.0n w=300n m=1
MMI8 VSS net11 VSS VSS nch_dnw l=690.0n w=300n m=1
MM_u2 net5 net11 VSS VSS nch_dnw l=60n w=300n m=1
MMI7 VSS net11 VSS VSS nch_dnw l=690.0n w=300n m=1
.ENDS

************************************************************************
* Library Name: CoRDIA_ADC_01
* Cell Name:    DECAP_UNIT
* View Name:    schematic
************************************************************************

.SUBCKT DECAP_UNIT VDD VSS
*.PININFO VDD:B VSS:B
XI0[77] VDD VSS / DCAP32
XI0[76] VDD VSS / DCAP32
XI0[75] VDD VSS / DCAP32
XI0[74] VDD VSS / DCAP32
XI0[73] VDD VSS / DCAP32
XI0[72] VDD VSS / DCAP32
XI0[71] VDD VSS / DCAP32
XI0[70] VDD VSS / DCAP32
XI0[69] VDD VSS / DCAP32
XI0[68] VDD VSS / DCAP32
XI0[67] VDD VSS / DCAP32
XI0[66] VDD VSS / DCAP32
XI0[65] VDD VSS / DCAP32
XI0[64] VDD VSS / DCAP32
XI0[63] VDD VSS / DCAP32
XI0[62] VDD VSS / DCAP32
XI0[61] VDD VSS / DCAP32
XI0[60] VDD VSS / DCAP32
XI0[59] VDD VSS / DCAP32
XI0[58] VDD VSS / DCAP32
XI0[57] VDD VSS / DCAP32
XI0[56] VDD VSS / DCAP32
XI0[55] VDD VSS / DCAP32
XI0[54] VDD VSS / DCAP32
XI0[53] VDD VSS / DCAP32
XI0[52] VDD VSS / DCAP32
XI0[51] VDD VSS / DCAP32
XI0[50] VDD VSS / DCAP32
XI0[49] VDD VSS / DCAP32
XI0[48] VDD VSS / DCAP32
XI0[47] VDD VSS / DCAP32
XI0[46] VDD VSS / DCAP32
XI0[45] VDD VSS / DCAP32
XI0[44] VDD VSS / DCAP32
XI0[43] VDD VSS / DCAP32
XI0[42] VDD VSS / DCAP32
XI0[41] VDD VSS / DCAP32
XI0[40] VDD VSS / DCAP32
XI0[39] VDD VSS / DCAP32
XI0[38] VDD VSS / DCAP32
XI0[37] VDD VSS / DCAP32
XI0[36] VDD VSS / DCAP32
XI0[35] VDD VSS / DCAP32
XI0[34] VDD VSS / DCAP32
XI0[33] VDD VSS / DCAP32
XI0[32] VDD VSS / DCAP32
XI0[31] VDD VSS / DCAP32
XI0[30] VDD VSS / DCAP32
XI0[29] VDD VSS / DCAP32
XI0[28] VDD VSS / DCAP32
XI0[27] VDD VSS / DCAP32
XI0[26] VDD VSS / DCAP32
XI0[25] VDD VSS / DCAP32
XI0[24] VDD VSS / DCAP32
XI0[23] VDD VSS / DCAP32
XI0[22] VDD VSS / DCAP32
XI0[21] VDD VSS / DCAP32
XI0[20] VDD VSS / DCAP32
XI0[19] VDD VSS / DCAP32
XI0[18] VDD VSS / DCAP32
XI0[17] VDD VSS / DCAP32
XI0[16] VDD VSS / DCAP32
XI0[15] VDD VSS / DCAP32
XI0[14] VDD VSS / DCAP32
XI0[13] VDD VSS / DCAP32
XI0[12] VDD VSS / DCAP32
XI0[11] VDD VSS / DCAP32
XI0[10] VDD VSS / DCAP32
XI0[9] VDD VSS / DCAP32
XI0[8] VDD VSS / DCAP32
XI0[7] VDD VSS / DCAP32
XI0[6] VDD VSS / DCAP32
XI0[5] VDD VSS / DCAP32
XI0[4] VDD VSS / DCAP32
XI0[3] VDD VSS / DCAP32
XI0[2] VDD VSS / DCAP32
XI0[1] VDD VSS / DCAP32
XI0[0] VDD VSS / DCAP32
XI1[25] VDD VSS / DCAP16
XI1[24] VDD VSS / DCAP16
XI1[23] VDD VSS / DCAP16
XI1[22] VDD VSS / DCAP16
XI1[21] VDD VSS / DCAP16
XI1[20] VDD VSS / DCAP16
XI1[19] VDD VSS / DCAP16
XI1[18] VDD VSS / DCAP16
XI1[17] VDD VSS / DCAP16
XI1[16] VDD VSS / DCAP16
XI1[15] VDD VSS / DCAP16
XI1[14] VDD VSS / DCAP16
XI1[13] VDD VSS / DCAP16
XI1[12] VDD VSS / DCAP16
XI1[11] VDD VSS / DCAP16
XI1[10] VDD VSS / DCAP16
XI1[9] VDD VSS / DCAP16
XI1[8] VDD VSS / DCAP16
XI1[7] VDD VSS / DCAP16
XI1[6] VDD VSS / DCAP16
XI1[5] VDD VSS / DCAP16
XI1[4] VDD VSS / DCAP16
XI1[3] VDD VSS / DCAP16
XI1[2] VDD VSS / DCAP16
XI1[1] VDD VSS / DCAP16
XI1[0] VDD VSS / DCAP16
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    TIEHLVT
* View Name:    schematic
************************************************************************

.SUBCKT TIEHLVT VDD VSS Z
*.PININFO Z:O VDD:B VSS:B
MM_u2 net7 net7 VSS VSS nch_lvt l=60n w=410.0n m=1
MM_u1 Z net7 VDD VDD pch_lvt l=60n w=540.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt_dnw
* Cell Name:    CKXOR2D4LVT_dnw
* View Name:    schematic
************************************************************************

.SUBCKT CKXOR2D4LVT_dnw A1 A2 VDD VSS Z
*.PININFO A1:I A2:I Z:O VDD:B VSS:B
MMM_u4_3-M_u3 Z net20 VDD VDD pch_lvt l=60n w=520.0n m=1
MMM_u2_1-M_u3 net97 A2 VDD VDD pch_lvt l=60n w=520.0n m=1
MMM_u2_0-M_u3 net97 A2 VDD VDD pch_lvt l=60n w=520.0n m=1
MMM_u2_2-M_u3 net97 A2 VDD VDD pch_lvt l=60n w=520.0n m=1
MMM_u5-M_u3 net61 net97 VDD VDD pch_lvt l=60n w=520.0n m=1
MMM_u6_0-M_u2 net97 A1 net20 VDD pch_lvt l=60n w=440.0n m=1
MMM_u4_1-M_u3 Z net20 VDD VDD pch_lvt l=60n w=520.0n m=1
MMM_u6_1-M_u2 net97 A1 net20 VDD pch_lvt l=60n w=440.0n m=1
MMM_u8-M_u3 net63 A1 VDD VDD pch_lvt l=60n w=520.0n m=1
MMM_u4_0-M_u3 Z net20 VDD VDD pch_lvt l=60n w=520.0n m=1
MMMI0_1-M_u2 net61 net63 net20 VDD pch_lvt l=60n w=395.00n m=1
MMMI0_0-M_u2 net61 net63 net20 VDD pch_lvt l=60n w=395.00n m=1
MMM_u4_2-M_u3 Z net20 VDD VDD pch_lvt l=60n w=520.0n m=1
MMM_u6_0-M_u3 net97 net63 net20 VSS nch_lvt_dnw l=60n w=275.00n m=1
MMMI0_0-M_u3 net61 A1 net20 VSS nch_lvt_dnw l=60n w=275.00n m=1
MMM_u8-M_u2 net63 A1 VSS VSS nch_lvt_dnw l=60n w=390.0n m=1
MMM_u2_1-M_u2 net97 A2 VSS VSS nch_lvt_dnw l=60n w=390.0n m=1
MMM_u4_1-M_u2 Z net20 VSS VSS nch_lvt_dnw l=60n w=390.0n m=1
MMM_u4_2-M_u2 Z net20 VSS VSS nch_lvt_dnw l=60n w=390.0n m=1
MMM_u6_1-M_u3 net97 net63 net20 VSS nch_lvt_dnw l=60n w=275.00n m=1
MMM_u5-M_u2 net61 net97 VSS VSS nch_lvt_dnw l=60n w=390.0n m=1
MMMI0_1-M_u3 net61 A1 net20 VSS nch_lvt_dnw l=60n w=275.00n m=1
MMM_u2_2-M_u2 net97 A2 VSS VSS nch_lvt_dnw l=60n w=390.0n m=1
MMM_u4_3-M_u2 Z net20 VSS VSS nch_lvt_dnw l=60n w=390.0n m=1
MMM_u4_0-M_u2 Z net20 VSS VSS nch_lvt_dnw l=60n w=390.0n m=1
MMM_u2_0-M_u2 net97 A2 VSS VSS nch_lvt_dnw l=60n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt_dnw
* Cell Name:    CKXOR2D2LVT_dnw
* View Name:    schematic
************************************************************************

.SUBCKT CKXOR2D2LVT_dnw A1 A2 VDD VSS Z
*.PININFO A1:I A2:I Z:O VDD:B VSS:B
MMM_u6-M_u2 net25 A1 net11 VDD pch_lvt l=60n w=290.0n m=1
MMM_u5-M_u3 net5 net25 VDD VDD pch_lvt l=60n w=290.0n m=1
MMM_u4_1-M_u3 Z net11 VDD VDD pch_lvt l=60n w=520.0n m=1
MMM_u8-M_u3 net13 A1 VDD VDD pch_lvt l=60n w=520.0n m=1
MMM_u4_0-M_u3 Z net11 VDD VDD pch_lvt l=60n w=520.0n m=1
MMMI0-M_u2 net5 net13 net11 VDD pch_lvt l=60n w=290.0n m=1
MMM_u2-M_u3 net25 A2 VDD VDD pch_lvt l=60n w=520.0n m=1
MMM_u6-M_u3 net25 net13 net11 VSS nch_lvt_dnw l=60n w=195.00n m=1
MMMI0-M_u3 net5 A1 net11 VSS nch_lvt_dnw l=60n w=195.00n m=1
MMM_u8-M_u2 net13 A1 VSS VSS nch_lvt_dnw l=60n w=195.00n m=1
MMM_u4_1-M_u2 Z net11 VSS VSS nch_lvt_dnw l=60n w=390.0n m=1
MMM_u2-M_u2 net25 A2 VSS VSS nch_lvt_dnw l=60n w=390.0n m=1
MMM_u5-M_u2 net5 net25 VSS VSS nch_lvt_dnw l=60n w=195.00n m=1
MMM_u4_0-M_u2 Z net11 VSS VSS nch_lvt_dnw l=60n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: frida
* Cell Name:    capdriver
* View Name:    schematic
************************************************************************

.SUBCKT capdriver dac_drive[15] dac_drive[14] dac_drive[13] dac_drive[12] 
+ dac_drive[11] dac_drive[10] dac_drive[9] dac_drive[8] dac_drive[7] 
+ dac_drive[6] dac_drive[5] dac_drive[4] dac_drive[3] dac_drive[2] 
+ dac_drive[1] dac_drive[0] dac_drive_invert dac_state[15] dac_state[14] 
+ dac_state[13] dac_state[12] dac_state[11] dac_state[10] dac_state[9] 
+ dac_state[8] dac_state[7] dac_state[6] dac_state[5] dac_state[4] 
+ dac_state[3] dac_state[2] dac_state[1] dac_state[0] vdd_dac vss_dac
*.PININFO dac_drive_invert:I dac_state[15]:I dac_state[14]:I dac_state[13]:I 
*.PININFO dac_state[12]:I dac_state[11]:I dac_state[10]:I dac_state[9]:I 
*.PININFO dac_state[8]:I dac_state[7]:I dac_state[6]:I dac_state[5]:I 
*.PININFO dac_state[4]:I dac_state[3]:I dac_state[2]:I dac_state[1]:I 
*.PININFO dac_state[0]:I dac_drive[15]:O dac_drive[14]:O dac_drive[13]:O 
*.PININFO dac_drive[12]:O dac_drive[11]:O dac_drive[10]:O dac_drive[9]:O 
*.PININFO dac_drive[8]:O dac_drive[7]:O dac_drive[6]:O dac_drive[5]:O 
*.PININFO dac_drive[4]:O dac_drive[3]:O dac_drive[2]:O dac_drive[1]:O 
*.PININFO dac_drive[0]:O vdd_dac:B vss_dac:B
XXxor15_0 dac_drive_invert dac_state[15] vdd_dac vss_dac dac_drive[15] / 
+ CKXOR2D4LVT_dnw
XXxor15_1 dac_drive_invert dac_state[15] vdd_dac vss_dac dac_drive[15] / 
+ CKXOR2D4LVT_dnw
XXxor14_0 dac_drive_invert dac_state[14] vdd_dac vss_dac dac_drive[14] / 
+ CKXOR2D4LVT_dnw
XXxor14_1 dac_drive_invert dac_state[14] vdd_dac vss_dac dac_drive[14] / 
+ CKXOR2D4LVT_dnw
XXxor13 dac_drive_invert dac_state[13] vdd_dac vss_dac dac_drive[13] / 
+ CKXOR2D4LVT_dnw
XXxor12 dac_drive_invert dac_state[12] vdd_dac vss_dac dac_drive[12] / 
+ CKXOR2D4LVT_dnw
XXxor11 dac_drive_invert dac_state[11] vdd_dac vss_dac dac_drive[11] / 
+ CKXOR2D2LVT_dnw
XXxor10 dac_drive_invert dac_state[10] vdd_dac vss_dac dac_drive[10] / 
+ CKXOR2D2LVT_dnw
XXxor9 dac_drive_invert dac_state[9] vdd_dac vss_dac dac_drive[9] / 
+ CKXOR2D2LVT_dnw
XXxor8 dac_drive_invert dac_state[8] vdd_dac vss_dac dac_drive[8] / 
+ CKXOR2D2LVT_dnw
XXxor7 dac_drive_invert dac_state[7] vdd_dac vss_dac dac_drive[7] / 
+ CKXOR2D2LVT_dnw
XXxor6 dac_drive_invert dac_state[6] vdd_dac vss_dac dac_drive[6] / 
+ CKXOR2D2LVT_dnw
XXxor5 dac_drive_invert dac_state[5] vdd_dac vss_dac dac_drive[5] / 
+ CKXOR2D2LVT_dnw
XXxor4 dac_drive_invert dac_state[4] vdd_dac vss_dac dac_drive[4] / 
+ CKXOR2D2LVT_dnw
XXxor3 dac_drive_invert dac_state[3] vdd_dac vss_dac dac_drive[3] / 
+ CKXOR2D2LVT_dnw
XXxor2 dac_drive_invert dac_state[2] vdd_dac vss_dac dac_drive[2] / 
+ CKXOR2D2LVT_dnw
XXxor1 dac_drive_invert dac_state[1] vdd_dac vss_dac dac_drive[1] / 
+ CKXOR2D2LVT_dnw
XXxor0 dac_drive_invert dac_state[0] vdd_dac vss_dac dac_drive[0] / 
+ CKXOR2D2LVT_dnw
.ENDS

************************************************************************
* Library Name: frida
* Cell Name:    caparray
* View Name:    schematic
************************************************************************

.SUBCKT caparray cap_botplate_diff[15] cap_botplate_diff[14] 
+ cap_botplate_diff[13] cap_botplate_diff[12] cap_botplate_diff[11] 
+ cap_botplate_diff[10] cap_botplate_diff[9] cap_botplate_diff[8] 
+ cap_botplate_diff[7] cap_botplate_diff[6] cap_botplate_diff[5] 
+ cap_botplate_diff[4] cap_botplate_diff[3] cap_botplate_diff[2] 
+ cap_botplate_diff[1] cap_botplate_diff[0] cap_botplate_main[15] 
+ cap_botplate_main[14] cap_botplate_main[13] cap_botplate_main[12] 
+ cap_botplate_main[11] cap_botplate_main[10] cap_botplate_main[9] 
+ cap_botplate_main[8] cap_botplate_main[7] cap_botplate_main[6] 
+ cap_botplate_main[5] cap_botplate_main[4] cap_botplate_main[3] 
+ cap_botplate_main[2] cap_botplate_main[1] cap_botplate_main[0] 
+ cap_shieldplate cap_topplate
*.PININFO cap_botplate_diff[15]:B cap_botplate_diff[14]:B 
*.PININFO cap_botplate_diff[13]:B cap_botplate_diff[12]:B 
*.PININFO cap_botplate_diff[11]:B cap_botplate_diff[10]:B 
*.PININFO cap_botplate_diff[9]:B cap_botplate_diff[8]:B cap_botplate_diff[7]:B 
*.PININFO cap_botplate_diff[6]:B cap_botplate_diff[5]:B cap_botplate_diff[4]:B 
*.PININFO cap_botplate_diff[3]:B cap_botplate_diff[2]:B cap_botplate_diff[1]:B 
*.PININFO cap_botplate_diff[0]:B cap_botplate_main[15]:B 
*.PININFO cap_botplate_main[14]:B cap_botplate_main[13]:B 
*.PININFO cap_botplate_main[12]:B cap_botplate_main[11]:B 
*.PININFO cap_botplate_main[10]:B cap_botplate_main[9]:B 
*.PININFO cap_botplate_main[8]:B cap_botplate_main[7]:B cap_botplate_main[6]:B 
*.PININFO cap_botplate_main[5]:B cap_botplate_main[4]:B cap_botplate_main[3]:B 
*.PININFO cap_botplate_main[2]:B cap_botplate_main[1]:B cap_botplate_main[0]:B 
*.PININFO cap_shieldplate:B cap_topplate:B

* Main and Diff capacitors based on exact weight calculations
* Weight 768: 768/64 = 12, so 12*0.4*(65+64) = 619.2f main, 12*0.4*(65-64) = 4.8f diff
Cmain15 cap_topplate cap_botplate_main[15] capacitor c=619.2f
Cdiff15 cap_topplate cap_botplate_diff[15] capacitor c=4.8f

* Weight 512: 512/64 = 8, so 8*0.4*(65+64) = 412.8f main, 8*0.4*(65-64) = 3.2f diff
Cmain14 cap_topplate cap_botplate_main[14] capacitor c=412.8f
Cdiff14 cap_topplate cap_botplate_diff[14] capacitor c=3.2f

* Weight 320: 320/64 = 5, so 5*0.4*(65+64) = 258f main, 5*0.4*(65-64) = 2f diff
Cmain13 cap_topplate cap_botplate_main[13] capacitor c=258f
Cdiff13 cap_topplate cap_botplate_diff[13] capacitor c=2f

* Weight 192: 192/64 = 3, so 3*0.4*(65+64) = 154.8f main, 3*0.4*(65-64) = 1.2f diff
Cmain12 cap_topplate cap_botplate_main[12] capacitor c=154.8f
Cdiff12 cap_topplate cap_botplate_diff[12] capacitor c=1.2f

* Weight 96: 64+32, so 0.4*(65+64)+0.4*(65+32) = 90.4f main, 0.4*(65-64)+0.4*(65-32) = 13.6f diff
Cmain11 cap_topplate cap_botplate_main[11] capacitor c=90.4f
Cdiff11 cap_topplate cap_botplate_diff[11] capacitor c=13.6f

* Weight 64: Single 64 section, 0.4*(65+64) = 51.6f main, 0.4*(65-64) = 0.4f diff
Cmain10 cap_topplate cap_botplate_main[10] capacitor c=51.6f
Cdiff10 cap_topplate cap_botplate_diff[10] capacitor c=0.4f

* Weight 32: 0.4*(65+32) = 38.8f main, 0.4*(65-32) = 13.2f diff
Cmain9 cap_topplate cap_botplate_main[9] capacitor c=38.8f
Cdiff9 cap_topplate cap_botplate_diff[9] capacitor c=13.2f

* Weight 24: 0.4*(65+24) = 35.6f main, 0.4*(65-24) = 16.4f diff
Cmain8 cap_topplate cap_botplate_main[8] capacitor c=35.6f
Cdiff8 cap_topplate cap_botplate_diff[8] capacitor c=16.4f

* Weight 12: 0.4*(65+12) = 30.8f main, 0.4*(65-12) = 21.2f diff
Cmain7 cap_topplate cap_botplate_main[7] capacitor c=30.8f
Cdiff7 cap_topplate cap_botplate_diff[7] capacitor c=21.2f

* Weight 10: 0.4*(65+10) = 30f main, 0.4*(65-10) = 22f diff
Cmain6 cap_topplate cap_botplate_main[6] capacitor c=30f
Cdiff6 cap_topplate cap_botplate_diff[6] capacitor c=22f

* Weight 5: 0.4*(65+5) = 28f main, 0.4*(65-5) = 24f diff
Cmain5 cap_topplate cap_botplate_main[5] capacitor c=28f
Cdiff5 cap_topplate cap_botplate_diff[5] capacitor c=24f

* Weight 4: 0.4*(65+4) = 27.6f main, 0.4*(65-4) = 24.4f diff
Cmain4 cap_topplate cap_botplate_main[4] capacitor c=27.6f
Cdiff4 cap_topplate cap_botplate_diff[4] capacitor c=24.4f

* Weight 4: Same as above
Cmain3 cap_topplate cap_botplate_main[3] capacitor c=27.6f
Cdiff3 cap_topplate cap_botplate_diff[3] capacitor c=24.4f

* Weight 2: 0.4*(65+2) = 26.8f main, 0.4*(65-2) = 25.2f diff
Cmain2 cap_topplate cap_botplate_main[2] capacitor c=26.8f
Cdiff2 cap_topplate cap_botplate_diff[2] capacitor c=25.2f

* Weight 1: 0.4*(65+1) = 26.4f main, 0.4*(65-1) = 25.6f diff
Cmain1 cap_topplate cap_botplate_main[1] capacitor c=26.4f
Cdiff1 cap_topplate cap_botplate_diff[1] capacitor c=25.6f

* Weight 1: Same as above
Cmain0 cap_topplate cap_botplate_main[0] capacitor c=26.4f
Cdiff0 cap_topplate cap_botplate_diff[0] capacitor c=25.6f

.ENDS

************************************************************************
* Library Name: frida
* Cell Name:    sampswitch
* View Name:    schematic
************************************************************************

.SUBCKT sampswitch clk clk_b vdd_a vin vout vss_a
*.PININFO clk:I clk_b:I vin:I vout:O vdd_a:B vss_a:B
MM1 vout clk_b vin vdd_a pch_lvt l=60n w=625.00n m=8
MM0 vout clk vin vss_a nch_lvt_dnw l=60n w=500n m=8
.ENDS

************************************************************************
* Library Name: tcbn65lp_dnw
* Cell Name:    NR2D2
* View Name:    schematic
************************************************************************

.SUBCKT NR2D2 A1 A2 VDD VSS ZN
*.PININFO A1:I A2:I ZN:O VDD:B VSS:B
MMI1_1-M_u2 ZN A1 net17 VDD pch l=60n w=530.0n m=1
MMI1_0-M_u1 net25 A2 VDD VDD pch l=60n w=530.0n m=1
MMI1_0-M_u2 ZN A1 net25 VDD pch l=60n w=530.0n m=1
MMI1_1-M_u1 net17 A2 VDD VDD pch l=60n w=530.0n m=1
MMI1_1-M_u3 ZN A2 VSS VSS nch_dnw l=60n w=390.0n m=1
MMI1_1-M_u4 ZN A1 VSS VSS nch_dnw l=60n w=390.0n m=1
MMI1_0-M_u4 ZN A1 VSS VSS nch_dnw l=60n w=390.0n m=1
MMI1_0-M_u3 ZN A2 VSS VSS nch_dnw l=60n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lp_dnw
* Cell Name:    CKND4
* View Name:    schematic
************************************************************************

.SUBCKT CKND4 I VDD VSS ZN
*.PININFO I:I ZN:O VDD:B VSS:B
MM_u2_1 ZN I VSS VSS nch_dnw l=60n w=310.0n m=1
MM_u2_3 ZN I VSS VSS nch_dnw l=60n w=310.0n m=1
MM_u2_0 ZN I VSS VSS nch_dnw l=60n w=310.0n m=1
MM_u2_2 ZN I VSS VSS nch_dnw l=60n w=310.0n m=1
MM_u1_0 ZN I VDD VDD pch l=60n w=520.0n m=1
MM_u1_3 ZN I VDD VDD pch l=60n w=520.0n m=1
MM_u1_2 ZN I VDD VDD pch l=60n w=520.0n m=1
MM_u1_1 ZN I VDD VDD pch l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lp_dnw
* Cell Name:    CKND8
* View Name:    schematic
************************************************************************

.SUBCKT CKND8 I VDD VSS ZN
*.PININFO I:I ZN:O VDD:B VSS:B
MM_u2_1 ZN I VSS VSS nch_dnw l=60n w=310.0n m=1
MM_u2_6 ZN I VSS VSS nch_dnw l=60n w=310.0n m=1
MM_u2_3 ZN I VSS VSS nch_dnw l=60n w=310.0n m=1
MM_u2_4 ZN I VSS VSS nch_dnw l=60n w=310.0n m=1
MM_u2_7 ZN I VSS VSS nch_dnw l=60n w=310.0n m=1
MM_u2_0 ZN I VSS VSS nch_dnw l=60n w=310.0n m=1
MM_u2_2 ZN I VSS VSS nch_dnw l=60n w=310.0n m=1
MM_u2_5 ZN I VSS VSS nch_dnw l=60n w=310.0n m=1
DDI3 VSS I ndio area=6.6e-14 pj=1.18e-06 m=1
MM_u1_7 ZN I VDD VDD pch l=60n w=520.0n m=1
MM_u1_0 ZN I VDD VDD pch l=60n w=520.0n m=1
MM_u1_3 ZN I VDD VDD pch l=60n w=520.0n m=1
MM_u1_2 ZN I VDD VDD pch l=60n w=520.0n m=1
MM_u1_4 ZN I VDD VDD pch l=60n w=520.0n m=1
MM_u1_6 ZN I VDD VDD pch l=60n w=520.0n m=1
MM_u1_1 ZN I VDD VDD pch l=60n w=520.0n m=1
MM_u1_5 ZN I VDD VDD pch l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: frida
* Cell Name:    comp_inverter_lvil
* View Name:    schematic
************************************************************************

.SUBCKT comp_inverter_lvil GND IN OUT VDD
*.PININFO IN:I OUT:O GND:B VDD:B
MMMN OUT IN GND GND nch_lvt_dnw l=60n w=390.0n m=1
MMMP OUT IN VDD VDD pch_hvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lp_dnw
* Cell Name:    DCAP8
* View Name:    schematic
************************************************************************

.SUBCKT DCAP8 VDD VSS
*.PININFO VDD:B VSS:B
MMI3 VDD net11 VDD VDD pch l=880.0n w=430.0n m=1
MM_u1 net9 net11 VDD VDD pch l=60n w=390.0n m=1
MMI4 VSS net9 VSS VSS nch_dnw l=880.0n w=300n m=1
MM_u2 net11 net9 VSS VSS nch_dnw l=60n w=300n m=1
.ENDS

************************************************************************
* Library Name: frida
* Cell Name:    comp_sr
* View Name:    schematic
************************************************************************

.SUBCKT comp_sr COMP_N COMP_P GND LATCH_N LATCH_P VDD
*.PININFO COMP_N:I COMP_P:I LATCH_N:O LATCH_P:O GND:B VDD:B
XXI30 net41 net38 VDD GND net35 / NR2D2
XXI31 net35 net42 VDD GND net38 / NR2D2
XXI45 net35 VDD GND net39 / CKND4
XXI48 net38 VDD GND net40 / CKND4
XXI46 net39 VDD GND LATCH_P / CKND8
XXI47 net40 VDD GND LATCH_N / CKND8
XXI22 GND COMP_P net41 VDD / comp_inverter_lvil
XXI0 GND COMP_N net42 VDD / comp_inverter_lvil
XXI1[5] VDD GND / DCAP8
XXI1[4] VDD GND / DCAP8
XXI1[3] VDD GND / DCAP8
XXI1[2] VDD GND / DCAP8
XXI1[1] VDD GND / DCAP8
XXI1[0] VDD GND / DCAP8
.ENDS

************************************************************************
* Library Name: frida
* Cell Name:    comp_latch
* View Name:    schematic
************************************************************************

.SUBCKT comp_latch CLK GND INN INP OUTN OUTP VDD
*.PININFO CLK:I INN:I INP:I OUTN:O OUTP:O GND:B VDD:B
MMM3 OUTN OUTP net031 GND nch_lvt_dnw l=350.0n w=750.0n m=4
MMM0 tail CLK GND GND nch_lvt_dnw l=800n w=550.0n m=1
MMM2 net037 INN tail GND nch_lvt_dnw l=300n w=1.1u m=4
MMM8[3] tail GND GND GND nch_lvt_dnw l=60n w=1.1u m=1
MMM8[2] tail GND GND GND nch_lvt_dnw l=60n w=1.1u m=1
MMM8[1] tail GND GND GND nch_lvt_dnw l=60n w=1.1u m=1
MMM8[0] tail GND GND GND nch_lvt_dnw l=60n w=1.1u m=1
MMM1 net031 INP tail GND nch_lvt_dnw l=300n w=1.1u m=4
MMM4 OUTP OUTN net037 GND nch_lvt_dnw l=350.0n w=750.0n m=4
MMS2 net037 CLK VDD VDD pch_lvt l=60n w=500n m=2
MMS4 OUTP CLK VDD VDD pch_lvt l=60n w=500n m=2
MMS1 net031 CLK VDD VDD pch_lvt l=60n w=500n m=2
MMM7 tail CLK VDD VDD pch_lvt l=60n w=500n m=1
MMM6 OUTP OUTN VDD VDD pch_lvt l=1u w=2u m=2
MMM5 OUTN OUTP VDD VDD pch_lvt l=1u w=2u m=2
MMS3 OUTN CLK VDD VDD pch_lvt l=60n w=500n m=2
.ENDS

************************************************************************
* Library Name: frida
* Cell Name:    comp
* View Name:    schematic
************************************************************************

.SUBCKT comp clk dout_n dout_p vdd_a vin_n vin_p vss_a
*.PININFO clk:I vin_n:I vin_p:I dout_n:O dout_p:O vdd_a:B vss_a:B
XXI3 COMP_N COMP_P vss_a dout_n dout_p vdd_a / comp_sr
XXLATCH clk vss_a vin_n vin_p COMP_N COMP_P vdd_a / comp_latch
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    BUFFD12LVT
* View Name:    schematic
************************************************************************

.SUBCKT BUFFD12LVT I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
MMU8_0-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_3-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_9-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_5-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_6-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u2_3-M_u2 net123 I VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u2_1-M_u2 net123 I VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_4-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_1-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u2_2-M_u2 net123 I VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_11-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u2_0-M_u2 net123 I VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_8-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_2-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_7-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_10-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_6-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_9-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_7-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_0-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2_1-M_u3 net123 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_4-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2_3-M_u3 net123 I VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2_0-M_u3 net123 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_11-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_8-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2_2-M_u3 net123 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_1-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_2-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_3-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_5-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_10-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    BUFFD0LVT
* View Name:    schematic
************************************************************************

.SUBCKT BUFFD0LVT I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
MMI2-M_u2 net5 I VSS VSS nch_lvt l=60n w=195.00n m=1
MMI1-M_u2 Z net5 VSS VSS nch_lvt l=60n w=195.00n m=1
MMI2-M_u3 net5 I VDD VDD pch_lvt l=60n w=260.0n m=1
MMI1-M_u3 Z net5 VDD VDD pch_lvt l=60n w=260.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    BUFFD2LVT
* View Name:    schematic
************************************************************************

.SUBCKT BUFFD2LVT I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
MM_u3_0-M_u3 Z net11 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_1-M_u3 Z net11 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2-M_u3 net11 I VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_1-M_u2 Z net11 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u2-M_u2 net11 I VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u3_0-M_u2 Z net11 VSS VSS nch_lvt l=60n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    CKBD2LVT
* View Name:    schematic
************************************************************************

.SUBCKT CKBD2LVT I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
MMU23_1 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MM_u15 net5 I VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_0 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MM_u3 net5 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_0 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_1 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    BUFFD4LVT
* View Name:    schematic
************************************************************************

.SUBCKT BUFFD4LVT I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
MM_u3_0-M_u3 Z net11 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2_1-M_u3 net11 I VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2_0-M_u3 net11 I VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_2-M_u3 Z net11 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_1-M_u3 Z net11 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_3-M_u3 Z net11 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_1-M_u2 Z net11 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u3_2-M_u2 Z net11 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u3_3-M_u2 Z net11 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u2_1-M_u2 net11 I VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u3_0-M_u2 Z net11 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u2_0-M_u2 net11 I VSS VSS nch_lvt l=60n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    DCAPLVT
* View Name:    schematic
************************************************************************

.SUBCKT DCAPLVT VDD VSS
*.PININFO VDD:B VSS:B
MM_u2 net7 net5 VSS VSS nch_lvt l=60n w=345.00n m=1
MM_u1 net5 net7 VDD VDD pch_lvt l=60n w=485.00n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    DCAP8LVT
* View Name:    schematic
************************************************************************

.SUBCKT DCAP8LVT VDD VSS
*.PININFO VDD:B VSS:B
MMI4 VSS net9 VSS VSS nch_lvt l=880.0n w=300n m=1
MM_u2 net11 net9 VSS VSS nch_lvt l=60n w=300n m=1
MMI3 VDD net11 VDD VDD pch_lvt l=880.0n w=430.0n m=1
MM_u1 net9 net11 VDD VDD pch_lvt l=60n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    DCAP4LVT
* View Name:    schematic
************************************************************************

.SUBCKT DCAP4LVT VDD VSS
*.PININFO VDD:B VSS:B
MMI4 VSS net9 VSS VSS nch_lvt l=80n w=330.0n m=1
MM_u2 net11 net9 VSS VSS nch_lvt l=60n w=330.0n m=1
MMI3 VDD net11 VDD VDD pch_lvt l=80n w=460.0n m=1
MM_u1 net9 net11 VDD VDD pch_lvt l=60n w=460.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    DCAP32LVT
* View Name:    schematic
************************************************************************

.SUBCKT DCAP32LVT VDD VSS
*.PININFO VDD:B VSS:B
MMI38 VSS net11 VSS VSS nch_lvt l=975.00n w=300n m=1
MMI6 VSS net11 VSS VSS nch_lvt l=975.00n w=300n m=1
MMI39 VSS net11 VSS VSS nch_lvt l=975.00n w=300n m=1
MMI37 VSS net11 VSS VSS nch_lvt l=975.00n w=300n m=1
MM_u2 net5 net11 VSS VSS nch_lvt l=60n w=300n m=1
MMI36 VSS net11 VSS VSS nch_lvt l=975.00n w=300n m=1
MMI33 VDD net5 VDD VDD pch_lvt l=975.00n w=430.0n m=1
MM_u1 net11 net5 VDD VDD pch_lvt l=60n w=390.0n m=1
MMI34 VDD net5 VDD VDD pch_lvt l=975.00n w=430.0n m=1
MMI35 VDD net5 VDD VDD pch_lvt l=975.00n w=430.0n m=1
MMI32 VDD net5 VDD VDD pch_lvt l=975.00n w=430.0n m=1
MMI26 VDD net5 VDD VDD pch_lvt l=975.00n w=430.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    INVD1LVT
* View Name:    schematic
************************************************************************

.SUBCKT INVD1LVT I VDD VSS ZN
*.PININFO I:I ZN:O VDD:B VSS:B
MMU1-M_u2 ZN I VSS VSS nch_lvt l=60n w=390.0n m=1
MMU1-M_u3 ZN I VDD VDD pch_lvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    CKLNQD1LVT
* View Name:    schematic
************************************************************************

.SUBCKT CKLNQD1LVT CP E Q TE VDD VSS
*.PININFO CP:I E:I TE:I Q:O VDD:B VSS:B
MMU19 net37 TE VSS VSS nch_lvt l=60n w=270.0n m=1
MMU20 net37 E VSS VSS nch_lvt l=60n w=270.0n m=1
MMI85-M_u4 net33 net63 VSS VSS nch_lvt l=60n w=215.00n m=1
MMI85-M_u3 net61 CP net33 VSS nch_lvt l=60n w=215.00n m=1
MMI82 net81 net9 net37 VSS nch_lvt l=60n w=270.0n m=1
MMU82-M_u2 net83 net9 VSS VSS nch_lvt l=60n w=195.00n m=1
MMI80-M_u2 net63 net81 VSS VSS nch_lvt l=60n w=215.00n m=1
MMI91 net13 net83 net81 VSS nch_lvt l=60n w=200n m=1
MMU81-M_u2 net9 CP VSS VSS nch_lvt l=60n w=195.00n m=1
MMI92 VSS net63 net13 VSS nch_lvt l=60n w=200n m=1
MMU75-M_u2 Q net61 VSS VSS nch_lvt l=60n w=215.00n m=1
MMU75-M_u3 Q net61 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU16 net81 net83 net45 VDD pch_lvt l=60n w=480.0n m=1
MMU82-M_u3 net83 net9 VDD VDD pch_lvt l=60n w=260.0n m=1
MMI85-M_u1 net61 CP VDD VDD pch_lvt l=60n w=350.0n m=1
MMU81-M_u3 net9 CP VDD VDD pch_lvt l=60n w=260.0n m=1
MMI81 net48 TE VDD VDD pch_lvt l=60n w=480.0n m=1
MMI85-M_u2 net61 net63 VDD VDD pch_lvt l=60n w=350.0n m=1
MMI80-M_u3 net63 net81 VDD VDD pch_lvt l=60n w=285.00n m=1
MMI90 net53 net9 net81 VDD pch_lvt l=60n w=200n m=1
MMI88 VDD net63 net53 VDD pch_lvt l=60n w=200n m=1
MMU17 net45 E net48 VDD pch_lvt l=60n w=480.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    CKND0LVT
* View Name:    schematic
************************************************************************

.SUBCKT CKND0LVT I VDD VSS ZN
*.PININFO I:I ZN:O VDD:B VSS:B
MM_u2 ZN I VSS VSS nch_lvt l=60n w=150.0n m=1
MM_u1 ZN I VDD VDD pch_lvt l=60n w=260.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    NR2D0LVT
* View Name:    schematic
************************************************************************

.SUBCKT NR2D0LVT A1 A2 VDD VSS ZN
*.PININFO A1:I A2:I ZN:O VDD:B VSS:B
MMI1-M_u3 ZN A2 VSS VSS nch_lvt l=60n w=195.00n m=1
MMI1-M_u4 ZN A1 VSS VSS nch_lvt l=60n w=195.00n m=1
MMI1-M_u1 net13 A2 VDD VDD pch_lvt l=60n w=260.0n m=1
MMI1-M_u2 ZN A1 net13 VDD pch_lvt l=60n w=260.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    CKND2D0LVT
* View Name:    schematic
************************************************************************

.SUBCKT CKND2D0LVT A1 A2 VDD VSS ZN
*.PININFO A1:I A2:I ZN:O VDD:B VSS:B
MMU1-M_u3 ZN A1 net1 VSS nch_lvt l=60n w=195.00n m=1
MMU1-M_u4 net1 A2 VSS VSS nch_lvt l=60n w=195.00n m=1
MMU1-M_u2 ZN A2 VDD VDD pch_lvt l=60n w=195.00n m=1
MMU1-M_u1 ZN A1 VDD VDD pch_lvt l=60n w=195.00n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    INVD2LVT
* View Name:    schematic
************************************************************************

.SUBCKT INVD2LVT I VDD VSS ZN
*.PININFO I:I ZN:O VDD:B VSS:B
MMU1_0-M_u2 ZN I VSS VSS nch_lvt l=60n w=390.0n m=1
MMU1_1-M_u2 ZN I VSS VSS nch_lvt l=60n w=390.0n m=1
MMU1_0-M_u3 ZN I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU1_1-M_u3 ZN I VDD VDD pch_lvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    ND2D2LVT
* View Name:    schematic
************************************************************************

.SUBCKT ND2D2LVT A1 A2 VDD VSS ZN
*.PININFO A1:I A2:I ZN:O VDD:B VSS:B
MMU3_1-M_u1 ZN A1 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU3_1-M_u2 ZN A2 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU3_0-M_u2 ZN A2 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU3_0-M_u1 ZN A1 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU3_0-M_u4 net20 A2 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU3_1-M_u3 ZN A1 net28 VSS nch_lvt l=60n w=390.0n m=1
MMU3_1-M_u4 net28 A2 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU3_0-M_u3 ZN A1 net20 VSS nch_lvt l=60n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    NR2D1LVT
* View Name:    schematic
************************************************************************

.SUBCKT NR2D1LVT A1 A2 VDD VSS ZN
*.PININFO A1:I A2:I ZN:O VDD:B VSS:B
MMI1-M_u3 ZN A2 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI1-M_u4 ZN A1 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI1-M_u1 net13 A2 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI1-M_u2 ZN A1 net13 VDD pch_lvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    INR2D2LVT
* View Name:    schematic
************************************************************************

.SUBCKT INR2D2LVT A1 B1 VDD VSS ZN
*.PININFO A1:I B1:I ZN:O VDD:B VSS:B
MMU1_0-M_u4 ZN B1 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU1_0-M_u3 ZN net5 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU1_1-M_u3 ZN net5 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU6-M_u2 net5 A1 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU1_1-M_u4 ZN B1 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU6-M_u3 net5 A1 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU1_0-M_u2 ZN B1 net36 VDD pch_lvt l=60n w=520.0n m=1
MMU1_0-M_u1 net36 net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU1_1-M_u1 net25 net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU1_1-M_u2 ZN B1 net25 VDD pch_lvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    IND2D0LVT
* View Name:    schematic
************************************************************************

.SUBCKT IND2D0LVT A1 B1 VDD VSS ZN
*.PININFO A1:I B1:I ZN:O VDD:B VSS:B
MMI2-M_u3 net9 A1 VDD VDD pch_lvt l=60n w=250.0n m=1
MMI11 VDD B1 ZN VDD pch_lvt l=60n w=250.0n m=1
MM_u16 VDD net9 ZN VDD pch_lvt l=60n w=250.0n m=1
MMI13 net21 net9 VSS VSS nch_lvt l=60n w=195.00n m=1
MMI2-M_u2 net9 A1 VSS VSS nch_lvt l=60n w=195.00n m=1
MMI12 ZN B1 net21 VSS nch_lvt l=60n w=195.00n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    NR2XD0LVT
* View Name:    schematic
************************************************************************

.SUBCKT NR2XD0LVT A1 A2 VDD VSS ZN
*.PININFO A1:I A2:I ZN:O VDD:B VSS:B
MMI1-M_u3 ZN A2 VSS VSS nch_lvt l=60n w=195.00n m=1
MMI1-M_u4 ZN A1 VSS VSS nch_lvt l=60n w=195.00n m=1
MMI1-M_u1 net13 A2 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI1-M_u2 ZN A1 net13 VDD pch_lvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    DFQD1LVT
* View Name:    schematic
************************************************************************

.SUBCKT DFQD1LVT CP D Q VDD VSS
*.PININFO CP:I D:I Q:O VDD:B VSS:B
MMI53-M_u2 net7 net13 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI4 net24 net63 VSS VSS nch_lvt l=60n w=370.0n m=1
MMI56 net37 net7 VSS VSS nch_lvt l=60n w=150.0n m=1
MMI13-M_u2 net11 net67 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI50 net11 net25 net13 VSS nch_lvt l=60n w=190.0n m=1
MMI32-M_u2 net25 net63 VSS VSS nch_lvt l=60n w=195.00n m=1
MMI5 net67 D net24 VSS nch_lvt l=60n w=370.0n m=1
MMI31-M_u2 net63 CP VSS VSS nch_lvt l=60n w=195.00n m=1
MMI49 net13 net63 net37 VSS nch_lvt l=60n w=150.0n m=1
MMI48 net9 net11 VSS VSS nch_lvt l=60n w=150.0n m=1
MMI27-M_u2 Q net7 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI47 net67 net25 net9 VSS nch_lvt l=60n w=150.0n m=1
MMI53-M_u3 net7 net13 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI32-M_u3 net25 net63 VDD VDD pch_lvt l=60n w=260.0n m=1
MMI43 net56 net11 VDD VDD pch_lvt l=60n w=150.0n m=1
MMI6 net67 D net49 VDD pch_lvt l=60n w=460.0n m=1
MMI31-M_u3 net63 CP VDD VDD pch_lvt l=60n w=260.0n m=1
MMI27-M_u3 Q net7 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI57 net13 net25 net72 VDD pch_lvt l=60n w=150.0n m=1
MMI13-M_u3 net11 net67 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI52 net11 net63 net13 VDD pch_lvt l=60n w=260.0n m=1
MMI51 net72 net7 VDD VDD pch_lvt l=60n w=150.0n m=1
MMI45 net67 net63 net56 VDD pch_lvt l=60n w=150.0n m=1
MMI7 net49 net25 VDD VDD pch_lvt l=60n w=460.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    EDFD2LVT
* View Name:    schematic
************************************************************************

.SUBCKT EDFD2LVT CP D E Q QN VDD VSS
*.PININFO CP:I D:I E:I Q:O QN:O VDD:B VSS:B
MMI75-M_u3 net51 net67 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI32-M_u3 net61 net11 VDD VDD pch_lvt l=60n w=260.0n m=1
MMI82-M_u3 net99 E VDD VDD pch_lvt l=60n w=290.0n m=1
MMI84 net93 D VDD VDD pch_lvt l=60n w=340.0n m=1
MMI29-M_u3 QN net51 VDD VDD pch_lvt l=60n w=1.04u m=1
MMI31-M_u3 net11 CP VDD VDD pch_lvt l=60n w=260.0n m=1
MMI27-M_u3 Q net67 VDD VDD pch_lvt l=60n w=1.04u m=1
MMI86 net5 E net33 VDD pch_lvt l=60n w=380.0n m=1
MMI85 net33 net51 VDD VDD pch_lvt l=60n w=380.0n m=1
MMI70 net29 net125 VDD VDD pch_lvt l=60n w=150.0n m=1
MMI73-M_u3 net67 net20 VDD VDD pch_lvt l=60n w=1.04u m=1
MMI67 net125 net11 net20 VDD pch_lvt l=60n w=340.0n m=1
MMI68 net51 net61 net20 VDD pch_lvt l=60n w=150.0n m=1
MMI74-M_u3 net125 net9 VDD VDD pch_lvt l=60n w=340.0n m=1
MMI69 net9 net11 net29 VDD pch_lvt l=60n w=150.0n m=1
MMI90 net5 net99 net93 VDD pch_lvt l=60n w=340.0n m=1
MMI83 net9 net61 net5 VDD pch_lvt l=60n w=340.0n m=1
MMI64 net72 net125 VSS VSS nch_lvt l=60n w=150.0n m=1
MMI29-M_u2 QN net51 VSS VSS nch_lvt l=60n w=780.0n m=1
MMI65 net125 net61 net20 VSS nch_lvt l=60n w=230.0n m=1
MMI82-M_u2 net99 E VSS VSS nch_lvt l=60n w=195.00n m=1
MMI89 net97 E net93 VSS nch_lvt l=60n w=210.0n m=1
MMI55 net51 net11 net20 VSS nch_lvt l=60n w=150.0n m=1
MMI77 net9 net11 net97 VSS nch_lvt l=60n w=290.0n m=1
MMI74-M_u2 net125 net9 VSS VSS nch_lvt l=60n w=150.0n m=1
MMI75-M_u2 net51 net67 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI81 net97 net99 net100 VSS nch_lvt l=60n w=350.0n m=1
MMI80 net93 D VSS VSS nch_lvt l=60n w=210.0n m=1
MMI32-M_u2 net61 net11 VSS VSS nch_lvt l=60n w=195.00n m=1
MMI31-M_u2 net11 CP VSS VSS nch_lvt l=60n w=195.00n m=1
MMI73-M_u2 net67 net20 VSS VSS nch_lvt l=60n w=780.0n m=1
MMI27-M_u2 Q net67 VSS VSS nch_lvt l=60n w=780.0n m=1
MMI78 net100 net51 VSS VSS nch_lvt l=60n w=350.0n m=1
MMI63 net9 net61 net72 VSS nch_lvt l=60n w=150.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    DCAP16LVT
* View Name:    schematic
************************************************************************

.SUBCKT DCAP16LVT VDD VSS
*.PININFO VDD:B VSS:B
MMI4 VSS net11 VSS VSS nch_lvt l=690.0n w=300n m=1
MMI8 VSS net11 VSS VSS nch_lvt l=690.0n w=300n m=1
MM_u2 net5 net11 VSS VSS nch_lvt l=60n w=300n m=1
MMI7 VSS net11 VSS VSS nch_lvt l=690.0n w=300n m=1
MMI3 VDD net5 VDD VDD pch_lvt l=690.0n w=430.0n m=1
MMI6 VDD net5 VDD VDD pch_lvt l=690.0n w=430.0n m=1
MM_u1 net11 net5 VDD VDD pch_lvt l=60n w=390.0n m=1
MMI5 VDD net5 VDD VDD pch_lvt l=690.0n w=430.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    DCAP64LVT
* View Name:    schematic
************************************************************************

.SUBCKT DCAP64LVT VDD VSS
*.PININFO VDD:B VSS:B
MMI54 VDD net11 VDD VDD pch_lvt l=915.00n w=430.0n m=1
MM_u1 net67 net11 VDD VDD pch_lvt l=60n w=390.0n m=1
MMI56 VDD net11 VDD VDD pch_lvt l=915.00n w=430.0n m=1
MMI55 VDD net11 VDD VDD pch_lvt l=915.00n w=430.0n m=1
MMI39 VDD net11 VDD VDD pch_lvt l=915.00n w=430.0n m=1
MMI57 VDD net11 VDD VDD pch_lvt l=915.00n w=430.0n m=1
MMI58 VDD net11 VDD VDD pch_lvt l=915.00n w=430.0n m=1
MMI59 VDD net11 VDD VDD pch_lvt l=915.00n w=430.0n m=1
MMI53 VDD net11 VDD VDD pch_lvt l=915.00n w=430.0n m=1
MMI50 VDD net11 VDD VDD pch_lvt l=915.00n w=430.0n m=1
MMI52 VDD net11 VDD VDD pch_lvt l=915.00n w=430.0n m=1
MMI51 VDD net11 VDD VDD pch_lvt l=915.00n w=430.0n m=1
MMI64 VSS net67 VSS VSS nch_lvt l=915.00n w=300n m=1
MMI65 VSS net67 VSS VSS nch_lvt l=915.00n w=300n m=1
MMI62 VSS net67 VSS VSS nch_lvt l=915.00n w=300n m=1
MMI67 VSS net67 VSS VSS nch_lvt l=915.00n w=300n m=1
MMI68 VSS net67 VSS VSS nch_lvt l=915.00n w=300n m=1
MMI60 VSS net67 VSS VSS nch_lvt l=915.00n w=300n m=1
MMI66 VSS net67 VSS VSS nch_lvt l=915.00n w=300n m=1
MMI69 VSS net67 VSS VSS nch_lvt l=915.00n w=300n m=1
MMI49 VSS net67 VSS VSS nch_lvt l=915.00n w=300n m=1
MMI61 VSS net67 VSS VSS nch_lvt l=915.00n w=300n m=1
MM_u2 net11 net67 VSS VSS nch_lvt l=60n w=300n m=1
MMI63 VSS net67 VSS VSS nch_lvt l=915.00n w=300n m=1
.ENDS

************************************************************************
* Library Name: frida
* Cell Name:    adc_digital
* View Name:    schematic
************************************************************************

.SUBCKT adc_digital clk_comp clk_samp_n clk_samp_n_b clk_samp_p clk_samp_p_b 
+ comp_out comp_out_n comp_out_p dac_astate_n[15] dac_astate_n[14] 
+ dac_astate_n[13] dac_astate_n[12] dac_astate_n[11] dac_astate_n[10] 
+ dac_astate_n[9] dac_astate_n[8] dac_astate_n[7] dac_astate_n[6] 
+ dac_astate_n[5] dac_astate_n[4] dac_astate_n[3] dac_astate_n[2] 
+ dac_astate_n[1] dac_astate_n[0] dac_astate_p[15] dac_astate_p[14] 
+ dac_astate_p[13] dac_astate_p[12] dac_astate_p[11] dac_astate_p[10] 
+ dac_astate_p[9] dac_astate_p[8] dac_astate_p[7] dac_astate_p[6] 
+ dac_astate_p[5] dac_astate_p[4] dac_astate_p[3] dac_astate_p[2] 
+ dac_astate_p[1] dac_astate_p[0] dac_bstate_n[15] dac_bstate_n[14] 
+ dac_bstate_n[13] dac_bstate_n[12] dac_bstate_n[11] dac_bstate_n[10] 
+ dac_bstate_n[9] dac_bstate_n[8] dac_bstate_n[7] dac_bstate_n[6] 
+ dac_bstate_n[5] dac_bstate_n[4] dac_bstate_n[3] dac_bstate_n[2] 
+ dac_bstate_n[1] dac_bstate_n[0] dac_bstate_p[15] dac_bstate_p[14] 
+ dac_bstate_p[13] dac_bstate_p[12] dac_bstate_p[11] dac_bstate_p[10] 
+ dac_bstate_p[9] dac_bstate_p[8] dac_bstate_p[7] dac_bstate_p[6] 
+ dac_bstate_p[5] dac_bstate_p[4] dac_bstate_p[3] dac_bstate_p[2] 
+ dac_bstate_p[1] dac_bstate_p[0] dac_diffcaps dac_invert_n_diff 
+ dac_invert_n_main dac_invert_p_diff dac_invert_p_main dac_mode 
+ dac_state_n_diff[15] dac_state_n_diff[14] dac_state_n_diff[13] 
+ dac_state_n_diff[12] dac_state_n_diff[11] dac_state_n_diff[10] 
+ dac_state_n_diff[9] dac_state_n_diff[8] dac_state_n_diff[7] 
+ dac_state_n_diff[6] dac_state_n_diff[5] dac_state_n_diff[4] 
+ dac_state_n_diff[3] dac_state_n_diff[2] dac_state_n_diff[1] 
+ dac_state_n_diff[0] dac_state_n_main[15] dac_state_n_main[14] 
+ dac_state_n_main[13] dac_state_n_main[12] dac_state_n_main[11] 
+ dac_state_n_main[10] dac_state_n_main[9] dac_state_n_main[8] 
+ dac_state_n_main[7] dac_state_n_main[6] dac_state_n_main[5] 
+ dac_state_n_main[4] dac_state_n_main[3] dac_state_n_main[2] 
+ dac_state_n_main[1] dac_state_n_main[0] dac_state_p_diff[15] 
+ dac_state_p_diff[14] dac_state_p_diff[13] dac_state_p_diff[12] 
+ dac_state_p_diff[11] dac_state_p_diff[10] dac_state_p_diff[9] 
+ dac_state_p_diff[8] dac_state_p_diff[7] dac_state_p_diff[6] 
+ dac_state_p_diff[5] dac_state_p_diff[4] dac_state_p_diff[3] 
+ dac_state_p_diff[2] dac_state_p_diff[1] dac_state_p_diff[0] 
+ dac_state_p_main[15] dac_state_p_main[14] dac_state_p_main[13] 
+ dac_state_p_main[12] dac_state_p_main[11] dac_state_p_main[10] 
+ dac_state_p_main[9] dac_state_p_main[8] dac_state_p_main[7] 
+ dac_state_p_main[6] dac_state_p_main[5] dac_state_p_main[4] 
+ dac_state_p_main[3] dac_state_p_main[2] dac_state_p_main[1] 
+ dac_state_p_main[0] en_comp en_init en_samp_n en_samp_p en_update seq_comp 
+ seq_init seq_samp seq_update vdd_d vss_d
*.PININFO comp_out_n:I comp_out_p:I dac_astate_n[15]:I dac_astate_n[14]:I 
*.PININFO dac_astate_n[13]:I dac_astate_n[12]:I dac_astate_n[11]:I 
*.PININFO dac_astate_n[10]:I dac_astate_n[9]:I dac_astate_n[8]:I 
*.PININFO dac_astate_n[7]:I dac_astate_n[6]:I dac_astate_n[5]:I 
*.PININFO dac_astate_n[4]:I dac_astate_n[3]:I dac_astate_n[2]:I 
*.PININFO dac_astate_n[1]:I dac_astate_n[0]:I dac_astate_p[15]:I 
*.PININFO dac_astate_p[14]:I dac_astate_p[13]:I dac_astate_p[12]:I 
*.PININFO dac_astate_p[11]:I dac_astate_p[10]:I dac_astate_p[9]:I 
*.PININFO dac_astate_p[8]:I dac_astate_p[7]:I dac_astate_p[6]:I 
*.PININFO dac_astate_p[5]:I dac_astate_p[4]:I dac_astate_p[3]:I 
*.PININFO dac_astate_p[2]:I dac_astate_p[1]:I dac_astate_p[0]:I 
*.PININFO dac_bstate_n[15]:I dac_bstate_n[14]:I dac_bstate_n[13]:I 
*.PININFO dac_bstate_n[12]:I dac_bstate_n[11]:I dac_bstate_n[10]:I 
*.PININFO dac_bstate_n[9]:I dac_bstate_n[8]:I dac_bstate_n[7]:I 
*.PININFO dac_bstate_n[6]:I dac_bstate_n[5]:I dac_bstate_n[4]:I 
*.PININFO dac_bstate_n[3]:I dac_bstate_n[2]:I dac_bstate_n[1]:I 
*.PININFO dac_bstate_n[0]:I dac_bstate_p[15]:I dac_bstate_p[14]:I 
*.PININFO dac_bstate_p[13]:I dac_bstate_p[12]:I dac_bstate_p[11]:I 
*.PININFO dac_bstate_p[10]:I dac_bstate_p[9]:I dac_bstate_p[8]:I 
*.PININFO dac_bstate_p[7]:I dac_bstate_p[6]:I dac_bstate_p[5]:I 
*.PININFO dac_bstate_p[4]:I dac_bstate_p[3]:I dac_bstate_p[2]:I 
*.PININFO dac_bstate_p[1]:I dac_bstate_p[0]:I dac_diffcaps:I dac_mode:I 
*.PININFO en_comp:I en_init:I en_samp_n:I en_samp_p:I en_update:I seq_comp:I 
*.PININFO seq_init:I seq_samp:I seq_update:I clk_comp:O clk_samp_n:O 
*.PININFO clk_samp_n_b:O clk_samp_p:O clk_samp_p_b:O comp_out:O 
*.PININFO dac_invert_n_diff:O dac_invert_n_main:O dac_invert_p_diff:O 
*.PININFO dac_invert_p_main:O dac_state_n_diff[15]:O dac_state_n_diff[14]:O 
*.PININFO dac_state_n_diff[13]:O dac_state_n_diff[12]:O dac_state_n_diff[11]:O 
*.PININFO dac_state_n_diff[10]:O dac_state_n_diff[9]:O dac_state_n_diff[8]:O 
*.PININFO dac_state_n_diff[7]:O dac_state_n_diff[6]:O dac_state_n_diff[5]:O 
*.PININFO dac_state_n_diff[4]:O dac_state_n_diff[3]:O dac_state_n_diff[2]:O 
*.PININFO dac_state_n_diff[1]:O dac_state_n_diff[0]:O dac_state_n_main[15]:O 
*.PININFO dac_state_n_main[14]:O dac_state_n_main[13]:O dac_state_n_main[12]:O 
*.PININFO dac_state_n_main[11]:O dac_state_n_main[10]:O dac_state_n_main[9]:O 
*.PININFO dac_state_n_main[8]:O dac_state_n_main[7]:O dac_state_n_main[6]:O 
*.PININFO dac_state_n_main[5]:O dac_state_n_main[4]:O dac_state_n_main[3]:O 
*.PININFO dac_state_n_main[2]:O dac_state_n_main[1]:O dac_state_n_main[0]:O 
*.PININFO dac_state_p_diff[15]:O dac_state_p_diff[14]:O dac_state_p_diff[13]:O 
*.PININFO dac_state_p_diff[12]:O dac_state_p_diff[11]:O dac_state_p_diff[10]:O 
*.PININFO dac_state_p_diff[9]:O dac_state_p_diff[8]:O dac_state_p_diff[7]:O 
*.PININFO dac_state_p_diff[6]:O dac_state_p_diff[5]:O dac_state_p_diff[4]:O 
*.PININFO dac_state_p_diff[3]:O dac_state_p_diff[2]:O dac_state_p_diff[1]:O 
*.PININFO dac_state_p_diff[0]:O dac_state_p_main[15]:O dac_state_p_main[14]:O 
*.PININFO dac_state_p_main[13]:O dac_state_p_main[12]:O dac_state_p_main[11]:O 
*.PININFO dac_state_p_main[10]:O dac_state_p_main[9]:O dac_state_p_main[8]:O 
*.PININFO dac_state_p_main[7]:O dac_state_p_main[6]:O dac_state_p_main[5]:O 
*.PININFO dac_state_p_main[4]:O dac_state_p_main[3]:O dac_state_p_main[2]:O 
*.PININFO dac_state_p_main[1]:O dac_state_p_main[0]:O vdd_d:B vss_d:B
XXclkgate_clkgate_comp_clkgate_cell_3 vdd_d vss_d net3 / TIELLVT
XX_04_1 vdd_d vss_d dac_invert_n_main / TIELLVT
XX_06_2 vdd_d vss_d dac_invert_p_main / TIELLVT
XXclkgate_clkgate_init_clkgate_cell_4 vdd_d vss_d net4 / TIELLVT
XXclkgate_clkgate_samp_n_clkgate_cell_5 vdd_d vss_d net5 / TIELLVT
XXclkgate_clkgate_samp_p_clkgate_cell_6 vdd_d vss_d net6 / TIELLVT
XXclkgate_clkgate_update_clkgate_cell_7 vdd_d vss_d net7 / TIELLVT
XXclkbuf_0_clk_update clk_update vdd_d vss_d clknet_0_clk_update / BUFFD12LVT
XXclkbuf_2_2_f_clk_update clknet_0_clk_update vdd_d vss_d 
+ clknet_2_2_leaf_clk_update / BUFFD12LVT
XXclkbuf_2_0_f_clk_update clknet_0_clk_update vdd_d vss_d 
+ clknet_2_0_leaf_clk_update / BUFFD12LVT
XXclkbuf_2_3_f_clk_update clknet_0_clk_update vdd_d vss_d 
+ clknet_2_3_leaf_clk_update / BUFFD12LVT
XXclkbuf_2_1_f_clk_update clknet_0_clk_update vdd_d vss_d 
+ clknet_2_1_leaf_clk_update / BUFFD12LVT
XX_03_ dac_diffcaps vdd_d vss_d net76 / BUFFD0LVT
XX_05_ dac_diffcaps vdd_d vss_d net77 / BUFFD0LVT
XXinput51 dac_bstate_n[3] vdd_d vss_d net51 / BUFFD2LVT
XXinput50 dac_bstate_n[2] vdd_d vss_d net50 / BUFFD2LVT
XXinput52 dac_bstate_n[4] vdd_d vss_d net52 / BUFFD2LVT
XXinput49 dac_bstate_n[1] vdd_d vss_d net49 / BUFFD2LVT
XXinput48 dac_bstate_n[15] vdd_d vss_d net48 / BUFFD2LVT
XXinput47 dac_bstate_n[14] vdd_d vss_d net47 / BUFFD2LVT
XXinput46 dac_bstate_n[13] vdd_d vss_d net46 / BUFFD2LVT
XXinput45 dac_bstate_n[12] vdd_d vss_d net45 / BUFFD2LVT
XXinput44 dac_bstate_n[11] vdd_d vss_d net44 / BUFFD2LVT
XXinput43 dac_bstate_n[10] vdd_d vss_d net43 / BUFFD2LVT
XXinput42 dac_bstate_n[0] vdd_d vss_d net42 / BUFFD2LVT
XXinput41 dac_astate_p[9] vdd_d vss_d net41 / BUFFD2LVT
XXinput40 dac_astate_p[8] vdd_d vss_d net40 / BUFFD2LVT
XXinput39 dac_astate_p[7] vdd_d vss_d net39 / BUFFD2LVT
XXinput38 dac_astate_p[6] vdd_d vss_d net38 / BUFFD2LVT
XXinput37 dac_astate_p[5] vdd_d vss_d net37 / BUFFD2LVT
XXinput36 dac_astate_p[4] vdd_d vss_d net36 / BUFFD2LVT
XXinput35 dac_astate_p[3] vdd_d vss_d net35 / BUFFD2LVT
XXinput34 dac_astate_p[2] vdd_d vss_d net34 / BUFFD2LVT
XXinput33 dac_astate_p[1] vdd_d vss_d net33 / BUFFD2LVT
XXinput32 dac_astate_p[15] vdd_d vss_d net32 / BUFFD2LVT
XXinput31 dac_astate_p[14] vdd_d vss_d net31 / BUFFD2LVT
XXinput30 dac_astate_p[13] vdd_d vss_d net30 / BUFFD2LVT
XXinput29 dac_astate_p[12] vdd_d vss_d net29 / BUFFD2LVT
XXinput28 dac_astate_p[11] vdd_d vss_d net28 / BUFFD2LVT
XXinput27 dac_astate_p[10] vdd_d vss_d net27 / BUFFD2LVT
XXinput26 dac_astate_p[0] vdd_d vss_d net26 / BUFFD2LVT
XXinput25 dac_astate_n[9] vdd_d vss_d net25 / BUFFD2LVT
XXinput24 dac_astate_n[8] vdd_d vss_d net24 / BUFFD2LVT
XXinput23 dac_astate_n[7] vdd_d vss_d net23 / BUFFD2LVT
XXinput22 dac_astate_n[6] vdd_d vss_d net22 / BUFFD2LVT
XXinput21 dac_astate_n[5] vdd_d vss_d net21 / BUFFD2LVT
XXinput20 dac_astate_n[4] vdd_d vss_d net20 / BUFFD2LVT
XXinput19 dac_astate_n[3] vdd_d vss_d net19 / BUFFD2LVT
XXinput18 dac_astate_n[2] vdd_d vss_d net18 / BUFFD2LVT
XXinput17 dac_astate_n[1] vdd_d vss_d net17 / BUFFD2LVT
XXinput16 dac_astate_n[15] vdd_d vss_d net16 / BUFFD2LVT
XXinput15 dac_astate_n[14] vdd_d vss_d net15 / BUFFD2LVT
XXinput14 dac_astate_n[13] vdd_d vss_d net14 / BUFFD2LVT
XXinput13 dac_astate_n[12] vdd_d vss_d net13 / BUFFD2LVT
XXinput12 dac_astate_n[11] vdd_d vss_d net12 / BUFFD2LVT
XXinput11 dac_astate_n[10] vdd_d vss_d net11 / BUFFD2LVT
XXinput10 dac_astate_n[0] vdd_d vss_d net10 / BUFFD2LVT
XXinput9 comp_out_p vdd_d vss_d net9 / BUFFD2LVT
XXinput8 comp_out_n vdd_d vss_d net8 / BUFFD2LVT
XXsampdriver_n_clk_buf_buf_cell clk_samp_n_raw vdd_d vss_d clk_samp_n / 
+ BUFFD2LVT
XXsampdriver_p_clk_buf_buf_cell clk_samp_p_raw vdd_d vss_d clk_samp_p / 
+ BUFFD2LVT
XXinput53 dac_bstate_n[5] vdd_d vss_d net53 / BUFFD2LVT
XXinput54 dac_bstate_n[6] vdd_d vss_d net54 / BUFFD2LVT
XXinput55 dac_bstate_n[7] vdd_d vss_d net55 / BUFFD2LVT
XXinput56 dac_bstate_n[8] vdd_d vss_d net56 / BUFFD2LVT
XXinput57 dac_bstate_n[9] vdd_d vss_d net57 / BUFFD2LVT
XXinput58 dac_bstate_p[0] vdd_d vss_d net58 / BUFFD2LVT
XXinput59 dac_bstate_p[10] vdd_d vss_d net59 / BUFFD2LVT
XXinput60 dac_bstate_p[11] vdd_d vss_d net60 / BUFFD2LVT
XXinput61 dac_bstate_p[12] vdd_d vss_d net61 / BUFFD2LVT
XXinput62 dac_bstate_p[13] vdd_d vss_d net62 / BUFFD2LVT
XXinput63 dac_bstate_p[14] vdd_d vss_d net63 / BUFFD2LVT
XXinput64 dac_bstate_p[15] vdd_d vss_d net64 / BUFFD2LVT
XXinput65 dac_bstate_p[1] vdd_d vss_d net65 / BUFFD2LVT
XXinput66 dac_bstate_p[2] vdd_d vss_d net66 / BUFFD2LVT
XXinput67 dac_bstate_p[3] vdd_d vss_d net67 / BUFFD2LVT
XXinput68 dac_bstate_p[4] vdd_d vss_d net68 / BUFFD2LVT
XXinput69 dac_bstate_p[5] vdd_d vss_d net69 / BUFFD2LVT
XXinput70 dac_bstate_p[6] vdd_d vss_d net70 / BUFFD2LVT
XXinput71 dac_bstate_p[7] vdd_d vss_d net71 / BUFFD2LVT
XXinput72 dac_bstate_p[8] vdd_d vss_d net72 / BUFFD2LVT
XXinput73 dac_bstate_p[9] vdd_d vss_d net73 / BUFFD2LVT
XXinput74 dac_mode vdd_d vss_d net74 / BUFFD2LVT
XXoutput75 net9 vdd_d vss_d comp_out / BUFFD2LVT
XXoutput76 net76 vdd_d vss_d dac_invert_n_diff / BUFFD2LVT
XXoutput77 net77 vdd_d vss_d dac_invert_p_diff / BUFFD2LVT
XXoutput78 net78 vdd_d vss_d dac_state_n_diff[0] / BUFFD2LVT
XXoutput79 net79 vdd_d vss_d dac_state_n_diff[10] / BUFFD2LVT
XXoutput80 net80 vdd_d vss_d dac_state_n_diff[11] / BUFFD2LVT
XXoutput81 net81 vdd_d vss_d dac_state_n_diff[12] / BUFFD2LVT
XXoutput82 net82 vdd_d vss_d dac_state_n_diff[13] / BUFFD2LVT
XXoutput83 net83 vdd_d vss_d dac_state_n_diff[14] / BUFFD2LVT
XXoutput84 net84 vdd_d vss_d dac_state_n_diff[15] / BUFFD2LVT
XXoutput85 net85 vdd_d vss_d dac_state_n_diff[1] / BUFFD2LVT
XXoutput86 net86 vdd_d vss_d dac_state_n_diff[2] / BUFFD2LVT
XXoutput87 net87 vdd_d vss_d dac_state_n_diff[3] / BUFFD2LVT
XXoutput88 net88 vdd_d vss_d dac_state_n_diff[4] / BUFFD2LVT
XXoutput89 net89 vdd_d vss_d dac_state_n_diff[5] / BUFFD2LVT
XXoutput90 net90 vdd_d vss_d dac_state_n_diff[6] / BUFFD2LVT
XXoutput91 net91 vdd_d vss_d dac_state_n_diff[7] / BUFFD2LVT
XXoutput92 net92 vdd_d vss_d dac_state_n_diff[8] / BUFFD2LVT
XXoutput93 net93 vdd_d vss_d dac_state_n_diff[9] / BUFFD2LVT
XXoutput94 net78 vdd_d vss_d dac_state_n_main[0] / BUFFD2LVT
XXoutput95 net79 vdd_d vss_d dac_state_n_main[10] / BUFFD2LVT
XXoutput96 net80 vdd_d vss_d dac_state_n_main[11] / BUFFD2LVT
XXoutput97 net81 vdd_d vss_d dac_state_n_main[12] / BUFFD2LVT
XXoutput98 net82 vdd_d vss_d dac_state_n_main[13] / BUFFD2LVT
XXoutput99 net83 vdd_d vss_d dac_state_n_main[14] / BUFFD2LVT
XXoutput100 net84 vdd_d vss_d dac_state_n_main[15] / BUFFD2LVT
XXoutput101 net85 vdd_d vss_d dac_state_n_main[1] / BUFFD2LVT
XXoutput102 net86 vdd_d vss_d dac_state_n_main[2] / BUFFD2LVT
XXoutput103 net87 vdd_d vss_d dac_state_n_main[3] / BUFFD2LVT
XXoutput104 net88 vdd_d vss_d dac_state_n_main[4] / BUFFD2LVT
XXoutput105 net89 vdd_d vss_d dac_state_n_main[5] / BUFFD2LVT
XXoutput106 net90 vdd_d vss_d dac_state_n_main[6] / BUFFD2LVT
XXoutput107 net91 vdd_d vss_d dac_state_n_main[7] / BUFFD2LVT
XXoutput108 net92 vdd_d vss_d dac_state_n_main[8] / BUFFD2LVT
XXoutput109 net93 vdd_d vss_d dac_state_n_main[9] / BUFFD2LVT
XXoutput110 net148 vdd_d vss_d dac_state_p_diff[0] / BUFFD2LVT
XXoutput111 net111 vdd_d vss_d dac_state_p_diff[10] / BUFFD2LVT
XXoutput112 net112 vdd_d vss_d dac_state_p_diff[11] / BUFFD2LVT
XXoutput113 net113 vdd_d vss_d dac_state_p_diff[12] / BUFFD2LVT
XXoutput114 net114 vdd_d vss_d dac_state_p_diff[13] / BUFFD2LVT
XXoutput115 net115 vdd_d vss_d dac_state_p_diff[14] / BUFFD2LVT
XXoutput116 net116 vdd_d vss_d dac_state_p_diff[15] / BUFFD2LVT
XXoutput117 net117 vdd_d vss_d dac_state_p_diff[1] / BUFFD2LVT
XXoutput118 net118 vdd_d vss_d dac_state_p_diff[2] / BUFFD2LVT
XXoutput119 net119 vdd_d vss_d dac_state_p_diff[3] / BUFFD2LVT
XXoutput120 net120 vdd_d vss_d dac_state_p_diff[4] / BUFFD2LVT
XXoutput121 net121 vdd_d vss_d dac_state_p_diff[5] / BUFFD2LVT
XXoutput122 net122 vdd_d vss_d dac_state_p_diff[6] / BUFFD2LVT
XXoutput123 net123 vdd_d vss_d dac_state_p_diff[7] / BUFFD2LVT
XXoutput124 net124 vdd_d vss_d dac_state_p_diff[8] / BUFFD2LVT
XXoutput125 net125 vdd_d vss_d dac_state_p_diff[9] / BUFFD2LVT
XXoutput126 net148 vdd_d vss_d dac_state_p_main[0] / BUFFD2LVT
XXoutput127 net111 vdd_d vss_d dac_state_p_main[10] / BUFFD2LVT
XXoutput128 net112 vdd_d vss_d dac_state_p_main[11] / BUFFD2LVT
XXoutput129 net113 vdd_d vss_d dac_state_p_main[12] / BUFFD2LVT
XXoutput130 net114 vdd_d vss_d dac_state_p_main[13] / BUFFD2LVT
XXoutput131 net115 vdd_d vss_d dac_state_p_main[14] / BUFFD2LVT
XXoutput132 net116 vdd_d vss_d dac_state_p_main[15] / BUFFD2LVT
XXoutput133 net117 vdd_d vss_d dac_state_p_main[1] / BUFFD2LVT
XXoutput134 net118 vdd_d vss_d dac_state_p_main[2] / BUFFD2LVT
XXoutput135 net119 vdd_d vss_d dac_state_p_main[3] / BUFFD2LVT
XXoutput136 net120 vdd_d vss_d dac_state_p_main[4] / BUFFD2LVT
XXoutput137 net121 vdd_d vss_d dac_state_p_main[5] / BUFFD2LVT
XXoutput138 net122 vdd_d vss_d dac_state_p_main[6] / BUFFD2LVT
XXoutput139 net123 vdd_d vss_d dac_state_p_main[7] / BUFFD2LVT
XXoutput140 net124 vdd_d vss_d dac_state_p_main[8] / BUFFD2LVT
XXoutput141 net125 vdd_d vss_d dac_state_p_main[9] / BUFFD2LVT
XXplace152 clk_init vdd_d vss_d net152 / CKBD2LVT
XXplace145 salogic_dual_dac_ff_dac_state_n_ff_D[6] vdd_d vss_d net145 / 
+ CKBD2LVT
XXplace147 salogic_dual_dac_ff_dac_state_n_ff_D[4] vdd_d vss_d net147 / 
+ CKBD2LVT
XXplace149 salogic_dual_041_ vdd_d vss_d net149 / CKBD2LVT
XXplace151 salogic_dual_032_ vdd_d vss_d net151 / CKBD2LVT
XXplace154 net74 vdd_d vss_d net154 / CKBD2LVT
XXplace144 salogic_dual_dac_ff_dac_state_n_ff_D[7] vdd_d vss_d net144 / 
+ CKBD2LVT
XXplace146 salogic_dual_dac_ff_dac_state_n_ff_D[5] vdd_d vss_d net146 / 
+ CKBD2LVT
XXplace148 net110 vdd_d vss_d net148 / CKBD2LVT
XXplace150 salogic_dual_032_ vdd_d vss_d net150 / CKBD2LVT
XXplace153 net152 vdd_d vss_d net153 / CKBD2LVT
XXplace155 net74 vdd_d vss_d net155 / CKBD2LVT
XXclkload0 clknet_2_1_leaf_clk_update vdd_d vss_d _unconnected_0 / BUFFD4LVT
XXclkload2 clknet_2_3_leaf_clk_update vdd_d vss_d _unconnected_1 / BUFFD4LVT
XXFILLER_0_13 vdd_d vss_d / DCAPLVT
XXFILLER_0_273 vdd_d vss_d / DCAPLVT
XXFILLER_2_163 vdd_d vss_d / DCAPLVT
XXFILLER_2_281 vdd_d vss_d / DCAPLVT
XXFILLER_2_297 vdd_d vss_d / DCAPLVT
XXFILLER_3_8 vdd_d vss_d / DCAPLVT
XXFILLER_3_17 vdd_d vss_d / DCAPLVT
XXFILLER_3_109 vdd_d vss_d / DCAPLVT
XXFILLER_3_167 vdd_d vss_d / DCAPLVT
XXFILLER_3_188 vdd_d vss_d / DCAPLVT
XXFILLER_4_297 vdd_d vss_d / DCAPLVT
XXFILLER_5_72 vdd_d vss_d / DCAPLVT
XXFILLER_5_166 vdd_d vss_d / DCAPLVT
XXFILLER_5_279 vdd_d vss_d / DCAPLVT
XXFILLER_6_4 vdd_d vss_d / DCAPLVT
XXFILLER_6_123 vdd_d vss_d / DCAPLVT
XXFILLER_6_186 vdd_d vss_d / DCAPLVT
XXFILLER_6_211 vdd_d vss_d / DCAPLVT
XXFILLER_6_222 vdd_d vss_d / DCAPLVT
XXFILLER_7_8 vdd_d vss_d / DCAPLVT
XXFILLER_7_159 vdd_d vss_d / DCAPLVT
XXFILLER_7_268 vdd_d vss_d / DCAPLVT
XXFILLER_7_297 vdd_d vss_d / DCAPLVT
XXFILLER_8_74 vdd_d vss_d / DCAPLVT
XXFILLER_8_192 vdd_d vss_d / DCAPLVT
XXFILLER_8_254 vdd_d vss_d / DCAPLVT
XXFILLER_8_261 vdd_d vss_d / DCAPLVT
XXFILLER_10_12 vdd_d vss_d / DCAPLVT
XXFILLER_10_297 vdd_d vss_d / DCAPLVT
XXFILLER_11_44 vdd_d vss_d / DCAPLVT
XXFILLER_11_151 vdd_d vss_d / DCAPLVT
XXFILLER_11_186 vdd_d vss_d / DCAPLVT
XXFILLER_12_255 vdd_d vss_d / DCAPLVT
XXFILLER_12_277 vdd_d vss_d / DCAPLVT
XXFILLER_14_4 vdd_d vss_d / DCAPLVT
XXFILLER_14_36 vdd_d vss_d / DCAPLVT
XXFILLER_14_62 vdd_d vss_d / DCAPLVT
XXFILLER_14_157 vdd_d vss_d / DCAPLVT
XXFILLER_14_291 vdd_d vss_d / DCAPLVT
XXFILLER_15_28 vdd_d vss_d / DCAPLVT
XXFILLER_15_84 vdd_d vss_d / DCAPLVT
XXFILLER_15_277 vdd_d vss_d / DCAPLVT
XXFILLER_16_19 vdd_d vss_d / DCAPLVT
XXFILLER_16_217 vdd_d vss_d / DCAPLVT
XXFILLER_17_265 vdd_d vss_d / DCAPLVT
XXFILLER_17_280 vdd_d vss_d / DCAPLVT
XXFILLER_18_84 vdd_d vss_d / DCAPLVT
XXFILLER_19_0 vdd_d vss_d / DCAPLVT
XXFILLER_19_9 vdd_d vss_d / DCAPLVT
XXFILLER_19_57 vdd_d vss_d / DCAPLVT
XXFILLER_19_84 vdd_d vss_d / DCAPLVT
XXFILLER_20_40 vdd_d vss_d / DCAPLVT
XXFILLER_20_55 vdd_d vss_d / DCAPLVT
XXFILLER_20_261 vdd_d vss_d / DCAPLVT
XXFILLER_20_274 vdd_d vss_d / DCAPLVT
XXFILLER_21_45 vdd_d vss_d / DCAPLVT
XXFILLER_21_264 vdd_d vss_d / DCAPLVT
XXFILLER_22_273 vdd_d vss_d / DCAPLVT
XXFILLER_23_47 vdd_d vss_d / DCAPLVT
XXFILLER_23_256 vdd_d vss_d / DCAPLVT
XXFILLER_23_277 vdd_d vss_d / DCAPLVT
XXFILLER_24_44 vdd_d vss_d / DCAPLVT
XXFILLER_24_281 vdd_d vss_d / DCAPLVT
XXFILLER_25_246 vdd_d vss_d / DCAPLVT
XXFILLER_25_297 vdd_d vss_d / DCAPLVT
XXFILLER_26_26 vdd_d vss_d / DCAPLVT
XXFILLER_26_51 vdd_d vss_d / DCAPLVT
XXFILLER_0_103 vdd_d vss_d / DCAP8LVT
XXFILLER_0_215 vdd_d vss_d / DCAP8LVT
XXFILLER_1_0 vdd_d vss_d / DCAP8LVT
XXFILLER_1_226 vdd_d vss_d / DCAP8LVT
XXFILLER_1_286 vdd_d vss_d / DCAP8LVT
XXFILLER_2_0 vdd_d vss_d / DCAP8LVT
XXFILLER_2_155 vdd_d vss_d / DCAP8LVT
XXFILLER_2_223 vdd_d vss_d / DCAP8LVT
XXFILLER_2_243 vdd_d vss_d / DCAP8LVT
XXFILLER_3_0 vdd_d vss_d / DCAP8LVT
XXFILLER_3_40 vdd_d vss_d / DCAP8LVT
XXFILLER_3_101 vdd_d vss_d / DCAP8LVT
XXFILLER_3_155 vdd_d vss_d / DCAP8LVT
XXFILLER_3_180 vdd_d vss_d / DCAP8LVT
XXFILLER_3_232 vdd_d vss_d / DCAP8LVT
XXFILLER_4_124 vdd_d vss_d / DCAP8LVT
XXFILLER_4_151 vdd_d vss_d / DCAP8LVT
XXFILLER_4_260 vdd_d vss_d / DCAP8LVT
XXFILLER_4_273 vdd_d vss_d / DCAP8LVT
XXFILLER_4_289 vdd_d vss_d / DCAP8LVT
XXFILLER_5_31 vdd_d vss_d / DCAP8LVT
XXFILLER_5_60 vdd_d vss_d / DCAP8LVT
XXFILLER_5_214 vdd_d vss_d / DCAP8LVT
XXFILLER_5_257 vdd_d vss_d / DCAP8LVT
XXFILLER_5_292 vdd_d vss_d / DCAP8LVT
XXFILLER_6_80 vdd_d vss_d / DCAP8LVT
XXFILLER_6_203 vdd_d vss_d / DCAP8LVT
XXFILLER_6_245 vdd_d vss_d / DCAP8LVT
XXFILLER_7_0 vdd_d vss_d / DCAP8LVT
XXFILLER_8_37 vdd_d vss_d / DCAP8LVT
XXFILLER_8_56 vdd_d vss_d / DCAP8LVT
XXFILLER_8_170 vdd_d vss_d / DCAP8LVT
XXFILLER_8_246 vdd_d vss_d / DCAP8LVT
XXFILLER_9_49 vdd_d vss_d / DCAP8LVT
XXFILLER_9_116 vdd_d vss_d / DCAP8LVT
XXFILLER_10_0 vdd_d vss_d / DCAP8LVT
XXFILLER_10_35 vdd_d vss_d / DCAP8LVT
XXFILLER_10_48 vdd_d vss_d / DCAP8LVT
XXFILLER_10_289 vdd_d vss_d / DCAP8LVT
XXFILLER_11_0 vdd_d vss_d / DCAP8LVT
XXFILLER_11_36 vdd_d vss_d / DCAP8LVT
XXFILLER_12_0 vdd_d vss_d / DCAP8LVT
XXFILLER_12_139 vdd_d vss_d / DCAP8LVT
XXFILLER_13_129 vdd_d vss_d / DCAP8LVT
XXFILLER_13_235 vdd_d vss_d / DCAP8LVT
XXFILLER_13_253 vdd_d vss_d / DCAP8LVT
XXFILLER_14_20 vdd_d vss_d / DCAP8LVT
XXFILLER_14_43 vdd_d vss_d / DCAP8LVT
XXFILLER_14_267 vdd_d vss_d / DCAP8LVT
XXFILLER_15_35 vdd_d vss_d / DCAP8LVT
XXFILLER_15_217 vdd_d vss_d / DCAP8LVT
XXFILLER_15_254 vdd_d vss_d / DCAP8LVT
XXFILLER_17_0 vdd_d vss_d / DCAP8LVT
XXFILLER_17_73 vdd_d vss_d / DCAP8LVT
XXFILLER_17_272 vdd_d vss_d / DCAP8LVT
XXFILLER_17_286 vdd_d vss_d / DCAP8LVT
XXFILLER_18_0 vdd_d vss_d / DCAP8LVT
XXFILLER_18_72 vdd_d vss_d / DCAP8LVT
XXFILLER_19_45 vdd_d vss_d / DCAP8LVT
XXFILLER_19_258 vdd_d vss_d / DCAP8LVT
XXFILLER_20_32 vdd_d vss_d / DCAP8LVT
XXFILLER_20_47 vdd_d vss_d / DCAP8LVT
XXFILLER_21_13 vdd_d vss_d / DCAP8LVT
XXFILLER_21_33 vdd_d vss_d / DCAP8LVT
XXFILLER_21_77 vdd_d vss_d / DCAP8LVT
XXFILLER_23_244 vdd_d vss_d / DCAP8LVT
XXFILLER_23_265 vdd_d vss_d / DCAP8LVT
XXFILLER_23_286 vdd_d vss_d / DCAP8LVT
XXFILLER_24_32 vdd_d vss_d / DCAP8LVT
XXFILLER_24_53 vdd_d vss_d / DCAP8LVT
XXFILLER_24_238 vdd_d vss_d / DCAP8LVT
XXFILLER_24_257 vdd_d vss_d / DCAP8LVT
XXFILLER_24_290 vdd_d vss_d / DCAP8LVT
XXFILLER_25_7 vdd_d vss_d / DCAP8LVT
XXFILLER_25_23 vdd_d vss_d / DCAP8LVT
XXFILLER_25_43 vdd_d vss_d / DCAP8LVT
XXFILLER_26_0 vdd_d vss_d / DCAP8LVT
XXFILLER_26_292 vdd_d vss_d / DCAP8LVT
XXFILLER_0_136 vdd_d vss_d / DCAP4LVT
XXFILLER_0_111 vdd_d vss_d / DCAP4LVT
XXFILLER_0_223 vdd_d vss_d / DCAP4LVT
XXFILLER_0_238 vdd_d vss_d / DCAP4LVT
XXFILLER_0_261 vdd_d vss_d / DCAP4LVT
XXFILLER_0_294 vdd_d vss_d / DCAP4LVT
XXFILLER_1_8 vdd_d vss_d / DCAP4LVT
XXFILLER_1_20 vdd_d vss_d / DCAP4LVT
XXFILLER_1_32 vdd_d vss_d / DCAP4LVT
XXFILLER_1_44 vdd_d vss_d / DCAP4LVT
XXFILLER_1_110 vdd_d vss_d / DCAP4LVT
XXFILLER_1_137 vdd_d vss_d / DCAP4LVT
XXFILLER_1_258 vdd_d vss_d / DCAP4LVT
XXFILLER_1_294 vdd_d vss_d / DCAP4LVT
XXFILLER_2_32 vdd_d vss_d / DCAP4LVT
XXFILLER_2_172 vdd_d vss_d / DCAP4LVT
XXFILLER_2_231 vdd_d vss_d / DCAP4LVT
XXFILLER_2_265 vdd_d vss_d / DCAP4LVT
XXFILLER_2_277 vdd_d vss_d / DCAP4LVT
XXFILLER_3_48 vdd_d vss_d / DCAP4LVT
XXFILLER_3_141 vdd_d vss_d / DCAP4LVT
XXFILLER_3_163 vdd_d vss_d / DCAP4LVT
XXFILLER_4_0 vdd_d vss_d / DCAP4LVT
XXFILLER_4_40 vdd_d vss_d / DCAP4LVT
XXFILLER_4_52 vdd_d vss_d / DCAP4LVT
XXFILLER_4_188 vdd_d vss_d / DCAP4LVT
XXFILLER_5_7 vdd_d vss_d / DCAP4LVT
XXFILLER_5_19 vdd_d vss_d / DCAP4LVT
XXFILLER_5_68 vdd_d vss_d / DCAP4LVT
XXFILLER_5_188 vdd_d vss_d / DCAP4LVT
XXFILLER_5_265 vdd_d vss_d / DCAP4LVT
XXFILLER_5_275 vdd_d vss_d / DCAP4LVT
XXFILLER_6_0 vdd_d vss_d / DCAP4LVT
XXFILLER_6_13 vdd_d vss_d / DCAP4LVT
XXFILLER_6_68 vdd_d vss_d / DCAP4LVT
XXFILLER_6_146 vdd_d vss_d / DCAP4LVT
XXFILLER_6_218 vdd_d vss_d / DCAP4LVT
XXFILLER_6_296 vdd_d vss_d / DCAP4LVT
XXFILLER_7_155 vdd_d vss_d / DCAP4LVT
XXFILLER_7_283 vdd_d vss_d / DCAP4LVT
XXFILLER_7_293 vdd_d vss_d / DCAP4LVT
XXFILLER_8_0 vdd_d vss_d / DCAP4LVT
XXFILLER_8_70 vdd_d vss_d / DCAP4LVT
XXFILLER_8_106 vdd_d vss_d / DCAP4LVT
XXFILLER_8_118 vdd_d vss_d / DCAP4LVT
XXFILLER_8_184 vdd_d vss_d / DCAP4LVT
XXFILLER_8_284 vdd_d vss_d / DCAP4LVT
XXFILLER_8_296 vdd_d vss_d / DCAP4LVT
XXFILLER_9_0 vdd_d vss_d / DCAP4LVT
XXFILLER_9_124 vdd_d vss_d / DCAP4LVT
XXFILLER_9_161 vdd_d vss_d / DCAP4LVT
XXFILLER_9_194 vdd_d vss_d / DCAP4LVT
XXFILLER_9_256 vdd_d vss_d / DCAP4LVT
XXFILLER_9_281 vdd_d vss_d / DCAP4LVT
XXFILLER_10_8 vdd_d vss_d / DCAP4LVT
XXFILLER_10_56 vdd_d vss_d / DCAP4LVT
XXFILLER_10_114 vdd_d vss_d / DCAP4LVT
XXFILLER_10_197 vdd_d vss_d / DCAP4LVT
XXFILLER_10_275 vdd_d vss_d / DCAP4LVT
XXFILLER_11_8 vdd_d vss_d / DCAP4LVT
XXFILLER_11_112 vdd_d vss_d / DCAP4LVT
XXFILLER_11_182 vdd_d vss_d / DCAP4LVT
XXFILLER_11_263 vdd_d vss_d / DCAP4LVT
XXFILLER_12_30 vdd_d vss_d / DCAP4LVT
XXFILLER_12_74 vdd_d vss_d / DCAP4LVT
XXFILLER_12_170 vdd_d vss_d / DCAP4LVT
XXFILLER_12_241 vdd_d vss_d / DCAP4LVT
XXFILLER_12_273 vdd_d vss_d / DCAP4LVT
XXFILLER_12_290 vdd_d vss_d / DCAP4LVT
XXFILLER_13_0 vdd_d vss_d / DCAP4LVT
XXFILLER_13_137 vdd_d vss_d / DCAP4LVT
XXFILLER_13_174 vdd_d vss_d / DCAP4LVT
XXFILLER_13_243 vdd_d vss_d / DCAP4LVT
XXFILLER_13_280 vdd_d vss_d / DCAP4LVT
XXFILLER_13_287 vdd_d vss_d / DCAP4LVT
XXFILLER_14_0 vdd_d vss_d / DCAP4LVT
XXFILLER_14_92 vdd_d vss_d / DCAP4LVT
XXFILLER_14_126 vdd_d vss_d / DCAP4LVT
XXFILLER_14_170 vdd_d vss_d / DCAP4LVT
XXFILLER_14_259 vdd_d vss_d / DCAP4LVT
XXFILLER_14_281 vdd_d vss_d / DCAP4LVT
XXFILLER_15_16 vdd_d vss_d / DCAP4LVT
XXFILLER_15_24 vdd_d vss_d / DCAP4LVT
XXFILLER_15_80 vdd_d vss_d / DCAP4LVT
XXFILLER_15_273 vdd_d vss_d / DCAP4LVT
XXFILLER_16_0 vdd_d vss_d / DCAP4LVT
XXFILLER_16_83 vdd_d vss_d / DCAP4LVT
XXFILLER_16_213 vdd_d vss_d / DCAP4LVT
XXFILLER_16_265 vdd_d vss_d / DCAP4LVT
XXFILLER_16_290 vdd_d vss_d / DCAP4LVT
XXFILLER_17_81 vdd_d vss_d / DCAP4LVT
XXFILLER_17_261 vdd_d vss_d / DCAP4LVT
XXFILLER_17_294 vdd_d vss_d / DCAP4LVT
XXFILLER_18_8 vdd_d vss_d / DCAP4LVT
XXFILLER_18_80 vdd_d vss_d / DCAP4LVT
XXFILLER_18_213 vdd_d vss_d / DCAP4LVT
XXFILLER_18_268 vdd_d vss_d / DCAP4LVT
XXFILLER_19_53 vdd_d vss_d / DCAP4LVT
XXFILLER_19_80 vdd_d vss_d / DCAP4LVT
XXFILLER_19_266 vdd_d vss_d / DCAP4LVT
XXFILLER_19_280 vdd_d vss_d / DCAP4LVT
XXFILLER_19_290 vdd_d vss_d / DCAP4LVT
XXFILLER_20_0 vdd_d vss_d / DCAP4LVT
XXFILLER_20_245 vdd_d vss_d / DCAP4LVT
XXFILLER_20_290 vdd_d vss_d / DCAP4LVT
XXFILLER_21_0 vdd_d vss_d / DCAP4LVT
XXFILLER_21_21 vdd_d vss_d / DCAP4LVT
XXFILLER_21_41 vdd_d vss_d / DCAP4LVT
XXFILLER_21_229 vdd_d vss_d / DCAP4LVT
XXFILLER_21_249 vdd_d vss_d / DCAP4LVT
XXFILLER_21_294 vdd_d vss_d / DCAP4LVT
XXFILLER_22_0 vdd_d vss_d / DCAP4LVT
XXFILLER_22_51 vdd_d vss_d / DCAP4LVT
XXFILLER_22_269 vdd_d vss_d / DCAP4LVT
XXFILLER_23_0 vdd_d vss_d / DCAP4LVT
XXFILLER_23_19 vdd_d vss_d / DCAP4LVT
XXFILLER_23_56 vdd_d vss_d / DCAP4LVT
XXFILLER_23_252 vdd_d vss_d / DCAP4LVT
XXFILLER_23_273 vdd_d vss_d / DCAP4LVT
XXFILLER_23_294 vdd_d vss_d / DCAP4LVT
XXFILLER_24_40 vdd_d vss_d / DCAP4LVT
XXFILLER_24_246 vdd_d vss_d / DCAP4LVT
XXFILLER_24_265 vdd_d vss_d / DCAP4LVT
XXFILLER_24_277 vdd_d vss_d / DCAP4LVT
XXFILLER_25_31 vdd_d vss_d / DCAP4LVT
XXFILLER_25_242 vdd_d vss_d / DCAP4LVT
XXFILLER_25_261 vdd_d vss_d / DCAP4LVT
XXFILLER_26_47 vdd_d vss_d / DCAP4LVT
XXFILLER_26_260 vdd_d vss_d / DCAP4LVT
XXFILLER_26_270 vdd_d vss_d / DCAP4LVT
XXFILLER_26_282 vdd_d vss_d / DCAP4LVT
XXFILLER_0_183 vdd_d vss_d / DCAP32LVT
XXFILLER_0_71 vdd_d vss_d / DCAP32LVT
XXFILLER_1_62 vdd_d vss_d / DCAP32LVT
XXFILLER_2_66 vdd_d vss_d / DCAP32LVT
XXFILLER_4_76 vdd_d vss_d / DCAP32LVT
XXFILLER_7_53 vdd_d vss_d / DCAP32LVT
XXFILLER_7_123 vdd_d vss_d / DCAP32LVT
XXFILLER_7_215 vdd_d vss_d / DCAP32LVT
XXFILLER_8_214 vdd_d vss_d / DCAP32LVT
XXFILLER_9_84 vdd_d vss_d / DCAP32LVT
XXFILLER_10_66 vdd_d vss_d / DCAP32LVT
XXFILLER_10_149 vdd_d vss_d / DCAP32LVT
XXFILLER_11_80 vdd_d vss_d / DCAP32LVT
XXFILLER_12_107 vdd_d vss_d / DCAP32LVT
XXFILLER_12_209 vdd_d vss_d / DCAP32LVT
XXFILLER_13_33 vdd_d vss_d / DCAP32LVT
XXFILLER_14_227 vdd_d vss_d / DCAP32LVT
XXFILLER_16_35 vdd_d vss_d / DCAP32LVT
XXFILLER_17_213 vdd_d vss_d / DCAP32LVT
XXFILLER_20_213 vdd_d vss_d / DCAP32LVT
XXFILLER_22_237 vdd_d vss_d / DCAP32LVT
XXFILLER_24_0 vdd_d vss_d / DCAP32LVT
XXclkload1 clknet_2_2_leaf_clk_update vdd_d vss_d _unconnected_2 / INVD1LVT
XXclkgate_clkgate_comp_clkgate_cell seq_comp en_comp clk_comp net3 vdd_d vss_d 
+ / CKLNQD1LVT
XXclkgate_clkgate_init_clkgate_cell seq_init en_init clk_init net4 vdd_d vss_d 
+ / CKLNQD1LVT
XXclkgate_clkgate_samp_n_clkgate_cell seq_samp en_samp_n clk_samp_n_raw net5 
+ vdd_d vss_d / CKLNQD1LVT
XXclkgate_clkgate_samp_p_clkgate_cell seq_samp en_samp_p clk_samp_p_raw net6 
+ vdd_d vss_d / CKLNQD1LVT
XXclkgate_clkgate_update_clkgate_cell seq_update en_update clk_update net7 
+ vdd_d vss_d / CKLNQD1LVT
XXsalogic_dual_174_ salogic_dual_dac_cycle[1] vdd_d vss_d salogic_dual_015_ / 
+ CKND0LVT
XXsalogic_dual_177_ salogic_dual_dac_cycle[11] vdd_d vss_d salogic_dual_017_ / 
+ CKND0LVT
XXsalogic_dual_179_ salogic_dual_dac_cycle[12] vdd_d vss_d salogic_dual_018_ / 
+ CKND0LVT
XXsalogic_dual_181_ salogic_dual_dac_cycle[13] vdd_d vss_d salogic_dual_019_ / 
+ CKND0LVT
XXsalogic_dual_183_ salogic_dual_dac_cycle[14] vdd_d vss_d salogic_dual_020_ / 
+ CKND0LVT
XXsalogic_dual_185_ salogic_dual_dac_cycle[15] vdd_d vss_d salogic_dual_021_ / 
+ CKND0LVT
XXsalogic_dual_187_ salogic_dual_dac_cycle[2] vdd_d vss_d salogic_dual_022_ / 
+ CKND0LVT
XXsalogic_dual_189_ salogic_dual_dac_cycle[3] vdd_d vss_d salogic_dual_023_ / 
+ CKND0LVT
XXsalogic_dual_191_ salogic_dual_dac_cycle[4] vdd_d vss_d salogic_dual_024_ / 
+ CKND0LVT
XXsalogic_dual_193_ salogic_dual_dac_cycle[5] vdd_d vss_d salogic_dual_025_ / 
+ CKND0LVT
XXsalogic_dual_195_ salogic_dual_dac_cycle[6] vdd_d vss_d salogic_dual_026_ / 
+ CKND0LVT
XXsalogic_dual_197_ salogic_dual_dac_cycle[7] vdd_d vss_d salogic_dual_027_ / 
+ CKND0LVT
XXsalogic_dual_199_ salogic_dual_dac_cycle[8] vdd_d vss_d salogic_dual_028_ / 
+ CKND0LVT
XXsalogic_dual_201_ salogic_dual_dac_cycle[9] vdd_d vss_d salogic_dual_029_ / 
+ CKND0LVT
XXsalogic_dual_203_ salogic_dual_dac_cycle[10] vdd_d vss_d salogic_dual_030_ / 
+ CKND0LVT
XXsalogic_dual_209_ net42 vdd_d vss_d salogic_dual_035_ / CKND0LVT
XXsalogic_dual_222_ net58 vdd_d vss_d salogic_dual_046_ / CKND0LVT
XXsalogic_dual_227_ net43 vdd_d vss_d salogic_dual_050_ / CKND0LVT
XXsalogic_dual_233_ net59 vdd_d vss_d salogic_dual_054_ / CKND0LVT
XXsalogic_dual_238_ net44 vdd_d vss_d salogic_dual_058_ / CKND0LVT
XXsalogic_dual_244_ net60 vdd_d vss_d salogic_dual_062_ / CKND0LVT
XXsalogic_dual_249_ net45 vdd_d vss_d salogic_dual_066_ / CKND0LVT
XXsalogic_dual_255_ net61 vdd_d vss_d salogic_dual_070_ / CKND0LVT
XXsalogic_dual_260_ net46 vdd_d vss_d salogic_dual_074_ / CKND0LVT
XXsalogic_dual_266_ net62 vdd_d vss_d salogic_dual_078_ / CKND0LVT
XXsalogic_dual_271_ net47 vdd_d vss_d salogic_dual_082_ / CKND0LVT
XXsalogic_dual_279_ net63 vdd_d vss_d salogic_dual_088_ / CKND0LVT
XXsalogic_dual_284_ net48 vdd_d vss_d salogic_dual_092_ / CKND0LVT
XXsalogic_dual_290_ net64 vdd_d vss_d salogic_dual_096_ / CKND0LVT
XXsalogic_dual_295_ net49 vdd_d vss_d salogic_dual_100_ / CKND0LVT
XXsalogic_dual_301_ net65 vdd_d vss_d salogic_dual_104_ / CKND0LVT
XXsalogic_dual_306_ net50 vdd_d vss_d salogic_dual_108_ / CKND0LVT
XXsalogic_dual_312_ net66 vdd_d vss_d salogic_dual_112_ / CKND0LVT
XXsalogic_dual_317_ net51 vdd_d vss_d salogic_dual_116_ / CKND0LVT
XXsalogic_dual_323_ net67 vdd_d vss_d salogic_dual_120_ / CKND0LVT
XXsalogic_dual_328_ net52 vdd_d vss_d salogic_dual_124_ / CKND0LVT
XXsalogic_dual_336_ net68 vdd_d vss_d salogic_dual_130_ / CKND0LVT
XXsalogic_dual_341_ net53 vdd_d vss_d salogic_dual_134_ / CKND0LVT
XXsalogic_dual_347_ net69 vdd_d vss_d salogic_dual_138_ / CKND0LVT
XXsalogic_dual_352_ net54 vdd_d vss_d salogic_dual_142_ / CKND0LVT
XXsalogic_dual_358_ net70 vdd_d vss_d salogic_dual_146_ / CKND0LVT
XXsalogic_dual_363_ net55 vdd_d vss_d salogic_dual_150_ / CKND0LVT
XXsalogic_dual_369_ net71 vdd_d vss_d salogic_dual_154_ / CKND0LVT
XXsalogic_dual_374_ net56 vdd_d vss_d salogic_dual_158_ / CKND0LVT
XXsalogic_dual_380_ net72 vdd_d vss_d salogic_dual_162_ / CKND0LVT
XXsalogic_dual_385_ net57 vdd_d vss_d salogic_dual_166_ / CKND0LVT
XXsalogic_dual_391_ net73 vdd_d vss_d salogic_dual_170_ / CKND0LVT
XXsalogic_dual_176_ salogic_dual_015_ net152 vdd_d vss_d salogic_dual_000_ / 
+ NR2D0LVT
XXsalogic_dual_178_ salogic_dual_017_ net152 vdd_d vss_d salogic_dual_001_ / 
+ NR2D0LVT
XXsalogic_dual_180_ salogic_dual_018_ net152 vdd_d vss_d salogic_dual_002_ / 
+ NR2D0LVT
XXsalogic_dual_182_ salogic_dual_019_ net152 vdd_d vss_d salogic_dual_003_ / 
+ NR2D0LVT
XXsalogic_dual_184_ salogic_dual_020_ net153 vdd_d vss_d salogic_dual_004_ / 
+ NR2D0LVT
XXsalogic_dual_186_ salogic_dual_021_ net153 vdd_d vss_d salogic_dual_005_ / 
+ NR2D0LVT
XXsalogic_dual_188_ salogic_dual_022_ net152 vdd_d vss_d salogic_dual_006_ / 
+ NR2D0LVT
XXsalogic_dual_190_ salogic_dual_023_ net152 vdd_d vss_d salogic_dual_007_ / 
+ NR2D0LVT
XXsalogic_dual_192_ salogic_dual_024_ net153 vdd_d vss_d salogic_dual_008_ / 
+ NR2D0LVT
XXsalogic_dual_194_ salogic_dual_025_ net153 vdd_d vss_d salogic_dual_009_ / 
+ NR2D0LVT
XXsalogic_dual_196_ salogic_dual_026_ net153 vdd_d vss_d salogic_dual_010_ / 
+ NR2D0LVT
XXsalogic_dual_198_ salogic_dual_027_ net153 vdd_d vss_d salogic_dual_011_ / 
+ NR2D0LVT
XXsalogic_dual_200_ salogic_dual_028_ net152 vdd_d vss_d salogic_dual_012_ / 
+ NR2D0LVT
XXsalogic_dual_202_ salogic_dual_029_ net152 vdd_d vss_d salogic_dual_013_ / 
+ NR2D0LVT
XXsalogic_dual_204_ salogic_dual_030_ net152 vdd_d vss_d salogic_dual_014_ / 
+ NR2D0LVT
XXsalogic_dual_211_ salogic_dual_035_ net155 vdd_d vss_d salogic_dual_037_ / 
+ NR2D0LVT
XXsalogic_dual_214_ net150 net10 vdd_d vss_d salogic_dual_040_ / NR2D0LVT
XXsalogic_dual_223_ salogic_dual_046_ net154 vdd_d vss_d salogic_dual_047_ / 
+ NR2D0LVT
XXsalogic_dual_225_ net151 net26 vdd_d vss_d salogic_dual_049_ / NR2D0LVT
XXsalogic_dual_228_ salogic_dual_050_ net155 vdd_d vss_d salogic_dual_051_ / 
+ NR2D0LVT
XXsalogic_dual_230_ net150 net11 vdd_d vss_d salogic_dual_053_ / NR2D0LVT
XXsalogic_dual_234_ salogic_dual_054_ net154 vdd_d vss_d salogic_dual_055_ / 
+ NR2D0LVT
XXsalogic_dual_236_ net151 net27 vdd_d vss_d salogic_dual_057_ / NR2D0LVT
XXsalogic_dual_239_ salogic_dual_058_ net155 vdd_d vss_d salogic_dual_059_ / 
+ NR2D0LVT
XXsalogic_dual_241_ net150 net12 vdd_d vss_d salogic_dual_061_ / NR2D0LVT
XXsalogic_dual_245_ salogic_dual_062_ net154 vdd_d vss_d salogic_dual_063_ / 
+ NR2D0LVT
XXsalogic_dual_247_ net151 net28 vdd_d vss_d salogic_dual_065_ / NR2D0LVT
XXsalogic_dual_250_ salogic_dual_066_ net155 vdd_d vss_d salogic_dual_067_ / 
+ NR2D0LVT
XXsalogic_dual_252_ net150 net13 vdd_d vss_d salogic_dual_069_ / NR2D0LVT
XXsalogic_dual_256_ salogic_dual_070_ net154 vdd_d vss_d salogic_dual_071_ / 
+ NR2D0LVT
XXsalogic_dual_258_ net151 net29 vdd_d vss_d salogic_dual_073_ / NR2D0LVT
XXsalogic_dual_261_ salogic_dual_074_ net155 vdd_d vss_d salogic_dual_075_ / 
+ NR2D0LVT
XXsalogic_dual_263_ net150 net14 vdd_d vss_d salogic_dual_077_ / NR2D0LVT
XXsalogic_dual_267_ salogic_dual_078_ net154 vdd_d vss_d salogic_dual_079_ / 
+ NR2D0LVT
XXsalogic_dual_269_ net151 net30 vdd_d vss_d salogic_dual_081_ / NR2D0LVT
XXsalogic_dual_273_ salogic_dual_082_ net155 vdd_d vss_d salogic_dual_084_ / 
+ NR2D0LVT
XXsalogic_dual_280_ salogic_dual_088_ net154 vdd_d vss_d salogic_dual_089_ / 
+ NR2D0LVT
XXsalogic_dual_285_ salogic_dual_092_ net155 vdd_d vss_d salogic_dual_093_ / 
+ NR2D0LVT
XXsalogic_dual_291_ salogic_dual_096_ net154 vdd_d vss_d salogic_dual_097_ / 
+ NR2D0LVT
XXsalogic_dual_296_ salogic_dual_100_ net155 vdd_d vss_d salogic_dual_101_ / 
+ NR2D0LVT
XXsalogic_dual_302_ salogic_dual_104_ net154 vdd_d vss_d salogic_dual_105_ / 
+ NR2D0LVT
XXsalogic_dual_307_ salogic_dual_108_ net155 vdd_d vss_d salogic_dual_109_ / 
+ NR2D0LVT
XXsalogic_dual_313_ salogic_dual_112_ net154 vdd_d vss_d salogic_dual_113_ / 
+ NR2D0LVT
XXsalogic_dual_318_ salogic_dual_116_ net155 vdd_d vss_d salogic_dual_117_ / 
+ NR2D0LVT
XXsalogic_dual_324_ salogic_dual_120_ net154 vdd_d vss_d salogic_dual_121_ / 
+ NR2D0LVT
XXsalogic_dual_330_ salogic_dual_124_ net155 vdd_d vss_d salogic_dual_126_ / 
+ NR2D0LVT
XXsalogic_dual_331_ salogic_dual_033_ salogic_dual_126_ vdd_d vss_d 
+ salogic_dual_127_ / NR2D0LVT
XXsalogic_dual_333_ net150 net20 vdd_d vss_d salogic_dual_129_ / NR2D0LVT
XXsalogic_dual_334_ salogic_dual_127_ salogic_dual_129_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_D[4] / NR2D0LVT
XXsalogic_dual_337_ salogic_dual_130_ net154 vdd_d vss_d salogic_dual_131_ / 
+ NR2D0LVT
XXsalogic_dual_338_ salogic_dual_044_ salogic_dual_131_ vdd_d vss_d 
+ salogic_dual_132_ / NR2D0LVT
XXsalogic_dual_339_ net151 net36 vdd_d vss_d salogic_dual_133_ / NR2D0LVT
XXsalogic_dual_340_ salogic_dual_132_ salogic_dual_133_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_p_ff_D[4] / NR2D0LVT
XXsalogic_dual_342_ salogic_dual_134_ net155 vdd_d vss_d salogic_dual_135_ / 
+ NR2D0LVT
XXsalogic_dual_343_ salogic_dual_033_ salogic_dual_135_ vdd_d vss_d 
+ salogic_dual_136_ / NR2D0LVT
XXsalogic_dual_344_ net150 net21 vdd_d vss_d salogic_dual_137_ / NR2D0LVT
XXsalogic_dual_345_ salogic_dual_136_ salogic_dual_137_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_D[5] / NR2D0LVT
XXsalogic_dual_348_ salogic_dual_138_ net154 vdd_d vss_d salogic_dual_139_ / 
+ NR2D0LVT
XXsalogic_dual_349_ salogic_dual_044_ salogic_dual_139_ vdd_d vss_d 
+ salogic_dual_140_ / NR2D0LVT
XXsalogic_dual_350_ net151 net37 vdd_d vss_d salogic_dual_141_ / NR2D0LVT
XXsalogic_dual_351_ salogic_dual_140_ salogic_dual_141_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_p_ff_D[5] / NR2D0LVT
XXsalogic_dual_353_ salogic_dual_142_ net155 vdd_d vss_d salogic_dual_143_ / 
+ NR2D0LVT
XXsalogic_dual_354_ salogic_dual_033_ salogic_dual_143_ vdd_d vss_d 
+ salogic_dual_144_ / NR2D0LVT
XXsalogic_dual_355_ net150 net22 vdd_d vss_d salogic_dual_145_ / NR2D0LVT
XXsalogic_dual_356_ salogic_dual_144_ salogic_dual_145_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_D[6] / NR2D0LVT
XXsalogic_dual_359_ salogic_dual_146_ net154 vdd_d vss_d salogic_dual_147_ / 
+ NR2D0LVT
XXsalogic_dual_360_ salogic_dual_044_ salogic_dual_147_ vdd_d vss_d 
+ salogic_dual_148_ / NR2D0LVT
XXsalogic_dual_361_ net151 net38 vdd_d vss_d salogic_dual_149_ / NR2D0LVT
XXsalogic_dual_362_ salogic_dual_148_ salogic_dual_149_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_p_ff_D[6] / NR2D0LVT
XXsalogic_dual_364_ salogic_dual_150_ net155 vdd_d vss_d salogic_dual_151_ / 
+ NR2D0LVT
XXsalogic_dual_365_ salogic_dual_033_ salogic_dual_151_ vdd_d vss_d 
+ salogic_dual_152_ / NR2D0LVT
XXsalogic_dual_366_ net150 net23 vdd_d vss_d salogic_dual_153_ / NR2D0LVT
XXsalogic_dual_367_ salogic_dual_152_ salogic_dual_153_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_D[7] / NR2D0LVT
XXsalogic_dual_370_ salogic_dual_154_ net154 vdd_d vss_d salogic_dual_155_ / 
+ NR2D0LVT
XXsalogic_dual_371_ salogic_dual_044_ salogic_dual_155_ vdd_d vss_d 
+ salogic_dual_156_ / NR2D0LVT
XXsalogic_dual_372_ net151 net39 vdd_d vss_d salogic_dual_157_ / NR2D0LVT
XXsalogic_dual_373_ salogic_dual_156_ salogic_dual_157_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_p_ff_D[7] / NR2D0LVT
XXsalogic_dual_375_ salogic_dual_158_ net155 vdd_d vss_d salogic_dual_159_ / 
+ NR2D0LVT
XXsalogic_dual_376_ salogic_dual_033_ salogic_dual_159_ vdd_d vss_d 
+ salogic_dual_160_ / NR2D0LVT
XXsalogic_dual_377_ net150 net24 vdd_d vss_d salogic_dual_161_ / NR2D0LVT
XXsalogic_dual_378_ salogic_dual_160_ salogic_dual_161_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_D[8] / NR2D0LVT
XXsalogic_dual_381_ salogic_dual_162_ net154 vdd_d vss_d salogic_dual_163_ / 
+ NR2D0LVT
XXsalogic_dual_382_ salogic_dual_044_ salogic_dual_163_ vdd_d vss_d 
+ salogic_dual_164_ / NR2D0LVT
XXsalogic_dual_383_ net151 net40 vdd_d vss_d salogic_dual_165_ / NR2D0LVT
XXsalogic_dual_384_ salogic_dual_164_ salogic_dual_165_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_p_ff_D[8] / NR2D0LVT
XXsalogic_dual_386_ salogic_dual_166_ net155 vdd_d vss_d salogic_dual_167_ / 
+ NR2D0LVT
XXsalogic_dual_387_ salogic_dual_033_ salogic_dual_167_ vdd_d vss_d 
+ salogic_dual_168_ / NR2D0LVT
XXsalogic_dual_388_ net150 net25 vdd_d vss_d salogic_dual_169_ / NR2D0LVT
XXsalogic_dual_392_ salogic_dual_170_ net154 vdd_d vss_d salogic_dual_171_ / 
+ NR2D0LVT
XXsalogic_dual_389_ salogic_dual_168_ salogic_dual_169_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_D[9] / NR2D0LVT
XXsalogic_dual_393_ salogic_dual_044_ salogic_dual_171_ vdd_d vss_d 
+ salogic_dual_172_ / NR2D0LVT
XXsalogic_dual_394_ net151 net41 vdd_d vss_d salogic_dual_173_ / NR2D0LVT
XXsalogic_dual_395_ salogic_dual_172_ salogic_dual_173_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_p_ff_D[9] / NR2D0LVT
XXsalogic_dual_205_ net155 net9 vdd_d vss_d salogic_dual_031_ / CKND2D0LVT
XXsalogic_dual_219_ net8 net154 vdd_d vss_d salogic_dual_043_ / CKND2D0LVT
XXsalogic_dual_232_ salogic_dual_041_ salogic_dual_030_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_E[10] / CKND2D0LVT
XXsalogic_dual_243_ salogic_dual_041_ salogic_dual_017_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_E[11] / CKND2D0LVT
XXsalogic_dual_254_ salogic_dual_041_ salogic_dual_018_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_E[12] / CKND2D0LVT
XXsalogic_dual_265_ net149 salogic_dual_019_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_E[13] / CKND2D0LVT
XXsalogic_dual_278_ net149 salogic_dual_020_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_E[14] / CKND2D0LVT
XXsalogic_dual_289_ net149 salogic_dual_021_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_E[15] / CKND2D0LVT
XXsalogic_dual_300_ salogic_dual_041_ salogic_dual_015_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_E[1] / CKND2D0LVT
XXsalogic_dual_311_ net149 salogic_dual_022_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_E[2] / CKND2D0LVT
XXsalogic_dual_322_ net149 salogic_dual_023_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_E[3] / CKND2D0LVT
XXsalogic_dual_335_ net149 salogic_dual_024_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_E[4] / CKND2D0LVT
XXsalogic_dual_346_ net149 salogic_dual_025_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_E[5] / CKND2D0LVT
XXsalogic_dual_357_ net149 salogic_dual_026_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_E[6] / CKND2D0LVT
XXsalogic_dual_368_ net149 salogic_dual_027_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_E[7] / CKND2D0LVT
XXsalogic_dual_379_ net149 salogic_dual_028_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_E[8] / CKND2D0LVT
XXsalogic_dual_390_ salogic_dual_041_ salogic_dual_029_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_E[9] / CKND2D0LVT
XXsalogic_dual_206_ net153 vdd_d vss_d salogic_dual_032_ / INVD2LVT
XXsampdriver_n_clk_inv_inv_cell clk_samp_n_raw vdd_d vss_d clk_samp_n_b / 
+ INVD2LVT
XXsampdriver_p_clk_inv_inv_cell clk_samp_p_raw vdd_d vss_d clk_samp_p_b / 
+ INVD2LVT
XXsalogic_dual_207_ salogic_dual_031_ salogic_dual_032_ vdd_d vss_d 
+ salogic_dual_033_ / ND2D2LVT
XXsalogic_dual_220_ salogic_dual_043_ net151 vdd_d vss_d salogic_dual_044_ / 
+ ND2D2LVT
XXsalogic_dual_212_ salogic_dual_033_ salogic_dual_037_ vdd_d vss_d 
+ salogic_dual_038_ / NR2D1LVT
XXsalogic_dual_215_ salogic_dual_038_ salogic_dual_040_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_D[0] / NR2D1LVT
XXsalogic_dual_224_ salogic_dual_044_ salogic_dual_047_ vdd_d vss_d 
+ salogic_dual_048_ / NR2D1LVT
XXsalogic_dual_226_ salogic_dual_048_ salogic_dual_049_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_p_ff_D[0] / NR2D1LVT
XXsalogic_dual_229_ salogic_dual_033_ salogic_dual_051_ vdd_d vss_d 
+ salogic_dual_052_ / NR2D1LVT
XXsalogic_dual_231_ salogic_dual_052_ salogic_dual_053_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_D[10] / NR2D1LVT
XXsalogic_dual_235_ salogic_dual_044_ salogic_dual_055_ vdd_d vss_d 
+ salogic_dual_056_ / NR2D1LVT
XXsalogic_dual_237_ salogic_dual_056_ salogic_dual_057_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_p_ff_D[10] / NR2D1LVT
XXsalogic_dual_240_ salogic_dual_033_ salogic_dual_059_ vdd_d vss_d 
+ salogic_dual_060_ / NR2D1LVT
XXsalogic_dual_242_ salogic_dual_060_ salogic_dual_061_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_D[11] / NR2D1LVT
XXsalogic_dual_246_ salogic_dual_044_ salogic_dual_063_ vdd_d vss_d 
+ salogic_dual_064_ / NR2D1LVT
XXsalogic_dual_248_ salogic_dual_064_ salogic_dual_065_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_p_ff_D[11] / NR2D1LVT
XXsalogic_dual_251_ salogic_dual_033_ salogic_dual_067_ vdd_d vss_d 
+ salogic_dual_068_ / NR2D1LVT
XXsalogic_dual_253_ salogic_dual_068_ salogic_dual_069_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_D[12] / NR2D1LVT
XXsalogic_dual_257_ salogic_dual_044_ salogic_dual_071_ vdd_d vss_d 
+ salogic_dual_072_ / NR2D1LVT
XXsalogic_dual_259_ salogic_dual_072_ salogic_dual_073_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_p_ff_D[12] / NR2D1LVT
XXsalogic_dual_262_ salogic_dual_033_ salogic_dual_075_ vdd_d vss_d 
+ salogic_dual_076_ / NR2D1LVT
XXsalogic_dual_264_ salogic_dual_076_ salogic_dual_077_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_D[13] / NR2D1LVT
XXsalogic_dual_268_ salogic_dual_044_ salogic_dual_079_ vdd_d vss_d 
+ salogic_dual_080_ / NR2D1LVT
XXsalogic_dual_270_ salogic_dual_080_ salogic_dual_081_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_p_ff_D[13] / NR2D1LVT
XXsalogic_dual_274_ salogic_dual_033_ salogic_dual_084_ vdd_d vss_d 
+ salogic_dual_085_ / NR2D1LVT
XXsalogic_dual_277_ salogic_dual_085_ salogic_dual_087_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_D[14] / NR2D1LVT
XXsalogic_dual_281_ salogic_dual_044_ salogic_dual_089_ vdd_d vss_d 
+ salogic_dual_090_ / NR2D1LVT
XXsalogic_dual_283_ salogic_dual_090_ salogic_dual_091_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_p_ff_D[14] / NR2D1LVT
XXsalogic_dual_286_ salogic_dual_033_ salogic_dual_093_ vdd_d vss_d 
+ salogic_dual_094_ / NR2D1LVT
XXsalogic_dual_288_ salogic_dual_094_ salogic_dual_095_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_D[15] / NR2D1LVT
XXsalogic_dual_292_ salogic_dual_044_ salogic_dual_097_ vdd_d vss_d 
+ salogic_dual_098_ / NR2D1LVT
XXsalogic_dual_294_ salogic_dual_098_ salogic_dual_099_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_p_ff_D[15] / NR2D1LVT
XXsalogic_dual_297_ salogic_dual_033_ salogic_dual_101_ vdd_d vss_d 
+ salogic_dual_102_ / NR2D1LVT
XXsalogic_dual_299_ salogic_dual_102_ salogic_dual_103_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_D[1] / NR2D1LVT
XXsalogic_dual_303_ salogic_dual_044_ salogic_dual_105_ vdd_d vss_d 
+ salogic_dual_106_ / NR2D1LVT
XXsalogic_dual_305_ salogic_dual_106_ salogic_dual_107_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_p_ff_D[1] / NR2D1LVT
XXsalogic_dual_308_ salogic_dual_033_ salogic_dual_109_ vdd_d vss_d 
+ salogic_dual_110_ / NR2D1LVT
XXsalogic_dual_310_ salogic_dual_110_ salogic_dual_111_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_D[2] / NR2D1LVT
XXsalogic_dual_314_ salogic_dual_044_ salogic_dual_113_ vdd_d vss_d 
+ salogic_dual_114_ / NR2D1LVT
XXsalogic_dual_316_ salogic_dual_114_ salogic_dual_115_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_p_ff_D[2] / NR2D1LVT
XXsalogic_dual_319_ salogic_dual_033_ salogic_dual_117_ vdd_d vss_d 
+ salogic_dual_118_ / NR2D1LVT
XXsalogic_dual_321_ salogic_dual_118_ salogic_dual_119_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_D[3] / NR2D1LVT
XXsalogic_dual_325_ salogic_dual_044_ salogic_dual_121_ vdd_d vss_d 
+ salogic_dual_122_ / NR2D1LVT
XXsalogic_dual_327_ salogic_dual_122_ salogic_dual_123_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_p_ff_D[3] / NR2D1LVT
XXsalogic_dual_216_ net155 net152 vdd_d vss_d salogic_dual_041_ / INR2D2LVT
XXsalogic_dual_218_ salogic_dual_dac_cycle[0] salogic_dual_041_ vdd_d vss_d 
+ salogic_dual_dac_ff_dac_state_n_ff_E[0] / IND2D0LVT
XXsalogic_dual_276_ net150 net15 vdd_d vss_d salogic_dual_087_ / NR2XD0LVT
XXsalogic_dual_282_ net151 net31 vdd_d vss_d salogic_dual_091_ / NR2XD0LVT
XXsalogic_dual_287_ net150 net16 vdd_d vss_d salogic_dual_095_ / NR2XD0LVT
XXsalogic_dual_293_ net151 net32 vdd_d vss_d salogic_dual_099_ / NR2XD0LVT
XXsalogic_dual_298_ net150 net17 vdd_d vss_d salogic_dual_103_ / NR2XD0LVT
XXsalogic_dual_304_ net151 net33 vdd_d vss_d salogic_dual_107_ / NR2XD0LVT
XXsalogic_dual_309_ net150 net18 vdd_d vss_d salogic_dual_111_ / NR2XD0LVT
XXsalogic_dual_315_ net151 net34 vdd_d vss_d salogic_dual_115_ / NR2XD0LVT
XXsalogic_dual_320_ net150 net19 vdd_d vss_d salogic_dual_119_ / NR2XD0LVT
XXsalogic_dual_326_ net151 net35 vdd_d vss_d salogic_dual_123_ / NR2XD0LVT
X1 clknet_2_2_leaf_clk_update salogic_dual_000_ salogic_dual_dac_cycle[0] 
+ vdd_d vss_d / DFQD1LVT
X3 clknet_2_3_leaf_clk_update salogic_dual_001_ salogic_dual_dac_cycle[10] 
+ vdd_d vss_d / DFQD1LVT
X5 clknet_2_3_leaf_clk_update salogic_dual_002_ salogic_dual_dac_cycle[11] 
+ vdd_d vss_d / DFQD1LVT
X7 clknet_2_3_leaf_clk_update salogic_dual_003_ salogic_dual_dac_cycle[12] 
+ vdd_d vss_d / DFQD1LVT
X9 clknet_2_1_leaf_clk_update salogic_dual_004_ salogic_dual_dac_cycle[13] 
+ vdd_d vss_d / DFQD1LVT
X11 clknet_2_1_leaf_clk_update salogic_dual_005_ salogic_dual_dac_cycle[14] 
+ vdd_d vss_d / DFQD1LVT
X13 clknet_2_1_leaf_clk_update net153 salogic_dual_dac_cycle[15] vdd_d vss_d / 
+ DFQD1LVT
X15 clknet_2_2_leaf_clk_update salogic_dual_006_ salogic_dual_dac_cycle[1] 
+ vdd_d vss_d / DFQD1LVT
X17 clknet_2_0_leaf_clk_update salogic_dual_007_ salogic_dual_dac_cycle[2] 
+ vdd_d vss_d / DFQD1LVT
X19 clknet_2_0_leaf_clk_update salogic_dual_008_ salogic_dual_dac_cycle[3] 
+ vdd_d vss_d / DFQD1LVT
X21 clknet_2_0_leaf_clk_update salogic_dual_009_ salogic_dual_dac_cycle[4] 
+ vdd_d vss_d / DFQD1LVT
X23 clknet_2_0_leaf_clk_update salogic_dual_010_ salogic_dual_dac_cycle[5] 
+ vdd_d vss_d / DFQD1LVT
X25 clknet_2_0_leaf_clk_update salogic_dual_011_ salogic_dual_dac_cycle[6] 
+ vdd_d vss_d / DFQD1LVT
X27 clknet_2_1_leaf_clk_update salogic_dual_012_ salogic_dual_dac_cycle[7] 
+ vdd_d vss_d / DFQD1LVT
X29 clknet_2_0_leaf_clk_update salogic_dual_013_ salogic_dual_dac_cycle[8] 
+ vdd_d vss_d / DFQD1LVT
X31 clknet_2_2_leaf_clk_update salogic_dual_014_ salogic_dual_dac_cycle[9] 
+ vdd_d vss_d / DFQD1LVT
XXsalogic_dual_dac_ff_dac_state_n_ff_dffe[0] clknet_2_2_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_n_ff_D[0] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[0] net78 _unconnected_3 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_p_ff_dffe[0] clknet_2_2_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_p_ff_D[0] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[0] net110 _unconnected_4 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_n_ff_dffe[10] clknet_2_3_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_n_ff_D[10] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[10] net79 _unconnected_5 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_p_ff_dffe[10] clknet_2_3_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_p_ff_D[10] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[10] net111 _unconnected_6 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_n_ff_dffe[11] clknet_2_3_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_n_ff_D[11] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[11] net80 _unconnected_7 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_p_ff_dffe[11] clknet_2_3_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_p_ff_D[11] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[11] net112 _unconnected_8 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_n_ff_dffe[12] clknet_2_3_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_n_ff_D[12] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[12] net81 _unconnected_9 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_p_ff_dffe[12] clknet_2_3_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_p_ff_D[12] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[12] net113 _unconnected_10 vdd_d vss_d 
+ / EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_n_ff_dffe[13] clknet_2_3_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_n_ff_D[13] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[13] net82 _unconnected_11 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_p_ff_dffe[13] clknet_2_1_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_p_ff_D[13] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[13] net114 _unconnected_12 vdd_d vss_d 
+ / EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_n_ff_dffe[14] clknet_2_1_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_n_ff_D[14] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[14] net83 _unconnected_13 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_p_ff_dffe[14] clknet_2_1_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_p_ff_D[14] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[14] net115 _unconnected_14 vdd_d vss_d 
+ / EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_n_ff_dffe[15] clknet_2_1_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_n_ff_D[15] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[15] net84 _unconnected_15 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_p_ff_dffe[15] clknet_2_1_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_p_ff_D[15] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[15] net116 _unconnected_16 vdd_d vss_d 
+ / EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_n_ff_dffe[1] clknet_2_2_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_n_ff_D[1] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[1] net85 _unconnected_17 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_p_ff_dffe[1] clknet_2_2_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_p_ff_D[1] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[1] net117 _unconnected_18 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_n_ff_dffe[2] clknet_2_2_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_n_ff_D[2] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[2] net86 _unconnected_19 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_p_ff_dffe[2] clknet_2_0_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_p_ff_D[2] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[2] net118 _unconnected_20 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_n_ff_dffe[3] clknet_2_2_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_n_ff_D[3] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[3] net87 _unconnected_21 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_p_ff_dffe[3] clknet_2_0_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_p_ff_D[3] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[3] net119 _unconnected_22 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_n_ff_dffe[4] clknet_2_0_leaf_clk_update net147 
+ salogic_dual_dac_ff_dac_state_n_ff_E[4] net88 _unconnected_23 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_p_ff_dffe[4] clknet_2_0_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_p_ff_D[4] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[4] net120 _unconnected_24 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_n_ff_dffe[5] clknet_2_0_leaf_clk_update net146 
+ salogic_dual_dac_ff_dac_state_n_ff_E[5] net89 _unconnected_25 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_p_ff_dffe[5] clknet_2_0_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_p_ff_D[5] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[5] net121 _unconnected_26 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_n_ff_dffe[6] clknet_2_0_leaf_clk_update net145 
+ salogic_dual_dac_ff_dac_state_n_ff_E[6] net90 _unconnected_27 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_p_ff_dffe[6] clknet_2_0_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_p_ff_D[6] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[6] net122 _unconnected_28 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_n_ff_dffe[7] clknet_2_1_leaf_clk_update net144 
+ salogic_dual_dac_ff_dac_state_n_ff_E[7] net91 _unconnected_29 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_p_ff_dffe[7] clknet_2_1_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_p_ff_D[7] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[7] net123 _unconnected_30 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_n_ff_dffe[8] clknet_2_3_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_n_ff_D[8] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[8] net92 _unconnected_31 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_p_ff_dffe[8] clknet_2_2_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_p_ff_D[8] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[8] net124 _unconnected_32 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_n_ff_dffe[9] clknet_2_2_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_n_ff_D[9] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[9] net93 _unconnected_33 vdd_d vss_d / 
+ EDFD2LVT
XXsalogic_dual_dac_ff_dac_state_p_ff_dffe[9] clknet_2_2_leaf_clk_update 
+ salogic_dual_dac_ff_dac_state_p_ff_D[9] 
+ salogic_dual_dac_ff_dac_state_n_ff_E[9] net125 _unconnected_34 vdd_d vss_d / 
+ EDFD2LVT
XXFILLER_1_94 vdd_d vss_d / DCAP16LVT
XXFILLER_1_242 vdd_d vss_d / DCAP16LVT
XXFILLER_1_270 vdd_d vss_d / DCAP16LVT
XXFILLER_2_16 vdd_d vss_d / DCAP16LVT
XXFILLER_2_139 vdd_d vss_d / DCAP16LVT
XXFILLER_2_207 vdd_d vss_d / DCAP16LVT
XXFILLER_3_24 vdd_d vss_d / DCAP16LVT
XXFILLER_3_85 vdd_d vss_d / DCAP16LVT
XXFILLER_3_216 vdd_d vss_d / DCAP16LVT
XXFILLER_4_108 vdd_d vss_d / DCAP16LVT
XXFILLER_5_44 vdd_d vss_d / DCAP16LVT
XXFILLER_5_105 vdd_d vss_d / DCAP16LVT
XXFILLER_5_198 vdd_d vss_d / DCAP16LVT
XXFILLER_6_130 vdd_d vss_d / DCAP16LVT
XXFILLER_7_85 vdd_d vss_d / DCAP16LVT
XXFILLER_7_247 vdd_d vss_d / DCAP16LVT
XXFILLER_8_150 vdd_d vss_d / DCAP16LVT
XXFILLER_9_33 vdd_d vss_d / DCAP16LVT
XXFILLER_10_98 vdd_d vss_d / DCAP16LVT
XXFILLER_10_181 vdd_d vss_d / DCAP16LVT
XXFILLER_11_166 vdd_d vss_d / DCAP16LVT
XXFILLER_11_247 vdd_d vss_d / DCAP16LVT
XXFILLER_13_65 vdd_d vss_d / DCAP16LVT
XXFILLER_13_113 vdd_d vss_d / DCAP16LVT
XXFILLER_13_219 vdd_d vss_d / DCAP16LVT
XXFILLER_14_141 vdd_d vss_d / DCAP16LVT
XXFILLER_15_0 vdd_d vss_d / DCAP16LVT
XXFILLER_15_283 vdd_d vss_d / DCAP16LVT
XXFILLER_16_67 vdd_d vss_d / DCAP16LVT
XXFILLER_16_249 vdd_d vss_d / DCAP16LVT
XXFILLER_17_33 vdd_d vss_d / DCAP16LVT
XXFILLER_17_245 vdd_d vss_d / DCAP16LVT
XXFILLER_18_30 vdd_d vss_d / DCAP16LVT
XXFILLER_18_248 vdd_d vss_d / DCAP16LVT
XXFILLER_19_29 vdd_d vss_d / DCAP16LVT
XXFILLER_19_64 vdd_d vss_d / DCAP16LVT
XXFILLER_19_242 vdd_d vss_d / DCAP16LVT
XXFILLER_21_213 vdd_d vss_d / DCAP16LVT
XXFILLER_22_35 vdd_d vss_d / DCAP16LVT
XXFILLER_22_69 vdd_d vss_d / DCAP16LVT
XXFILLER_22_213 vdd_d vss_d / DCAP16LVT
XXFILLER_23_31 vdd_d vss_d / DCAP16LVT
XXFILLER_25_273 vdd_d vss_d / DCAP16LVT
XXFILLER_26_244 vdd_d vss_d / DCAP16LVT
XXFILLER_1_162 vdd_d vss_d / DCAP64LVT
XXFILLER_4_196 vdd_d vss_d / DCAP64LVT
XXFILLER_10_205 vdd_d vss_d / DCAP64LVT
.ENDS

************************************************************************
* Library Name: frida
* Cell Name:    adc
* View Name:    schematic
************************************************************************

.SUBCKT adc comp_out dac_astate_n[15] dac_astate_n[14] dac_astate_n[13] 
+ dac_astate_n[12] dac_astate_n[11] dac_astate_n[10] dac_astate_n[9] 
+ dac_astate_n[8] dac_astate_n[7] dac_astate_n[6] dac_astate_n[5] 
+ dac_astate_n[4] dac_astate_n[3] dac_astate_n[2] dac_astate_n[1] 
+ dac_astate_n[0] dac_astate_p[15] dac_astate_p[14] dac_astate_p[13] 
+ dac_astate_p[12] dac_astate_p[11] dac_astate_p[10] dac_astate_p[9] 
+ dac_astate_p[8] dac_astate_p[7] dac_astate_p[6] dac_astate_p[5] 
+ dac_astate_p[4] dac_astate_p[3] dac_astate_p[2] dac_astate_p[1] 
+ dac_astate_p[0] dac_bstate_n[15] dac_bstate_n[14] dac_bstate_n[13] 
+ dac_bstate_n[12] dac_bstate_n[11] dac_bstate_n[10] dac_bstate_n[9] 
+ dac_bstate_n[8] dac_bstate_n[7] dac_bstate_n[6] dac_bstate_n[5] 
+ dac_bstate_n[4] dac_bstate_n[3] dac_bstate_n[2] dac_bstate_n[1] 
+ dac_bstate_n[0] dac_bstate_p[15] dac_bstate_p[14] dac_bstate_p[13] 
+ dac_bstate_p[12] dac_bstate_p[11] dac_bstate_p[10] dac_bstate_p[9] 
+ dac_bstate_p[8] dac_bstate_p[7] dac_bstate_p[6] dac_bstate_p[5] 
+ dac_bstate_p[4] dac_bstate_p[3] dac_bstate_p[2] dac_bstate_p[1] 
+ dac_bstate_p[0] dac_diffcaps dac_mode en_comp en_init en_samp_n en_samp_p 
+ en_update seq_comp seq_init seq_samp seq_update vdd_a vdd_d vdd_dac vin_n 
+ vin_p vss_a vss_d vss_dac
*.PININFO dac_astate_n[15]:I dac_astate_n[14]:I dac_astate_n[13]:I 
*.PININFO dac_astate_n[12]:I dac_astate_n[11]:I dac_astate_n[10]:I 
*.PININFO dac_astate_n[9]:I dac_astate_n[8]:I dac_astate_n[7]:I 
*.PININFO dac_astate_n[6]:I dac_astate_n[5]:I dac_astate_n[4]:I 
*.PININFO dac_astate_n[3]:I dac_astate_n[2]:I dac_astate_n[1]:I 
*.PININFO dac_astate_n[0]:I dac_astate_p[15]:I dac_astate_p[14]:I 
*.PININFO dac_astate_p[13]:I dac_astate_p[12]:I dac_astate_p[11]:I 
*.PININFO dac_astate_p[10]:I dac_astate_p[9]:I dac_astate_p[8]:I 
*.PININFO dac_astate_p[7]:I dac_astate_p[6]:I dac_astate_p[5]:I 
*.PININFO dac_astate_p[4]:I dac_astate_p[3]:I dac_astate_p[2]:I 
*.PININFO dac_astate_p[1]:I dac_astate_p[0]:I dac_bstate_n[15]:I 
*.PININFO dac_bstate_n[14]:I dac_bstate_n[13]:I dac_bstate_n[12]:I 
*.PININFO dac_bstate_n[11]:I dac_bstate_n[10]:I dac_bstate_n[9]:I 
*.PININFO dac_bstate_n[8]:I dac_bstate_n[7]:I dac_bstate_n[6]:I 
*.PININFO dac_bstate_n[5]:I dac_bstate_n[4]:I dac_bstate_n[3]:I 
*.PININFO dac_bstate_n[2]:I dac_bstate_n[1]:I dac_bstate_n[0]:I 
*.PININFO dac_bstate_p[15]:I dac_bstate_p[14]:I dac_bstate_p[13]:I 
*.PININFO dac_bstate_p[12]:I dac_bstate_p[11]:I dac_bstate_p[10]:I 
*.PININFO dac_bstate_p[9]:I dac_bstate_p[8]:I dac_bstate_p[7]:I 
*.PININFO dac_bstate_p[6]:I dac_bstate_p[5]:I dac_bstate_p[4]:I 
*.PININFO dac_bstate_p[3]:I dac_bstate_p[2]:I dac_bstate_p[1]:I 
*.PININFO dac_bstate_p[0]:I dac_diffcaps:I dac_mode:I en_comp:I en_init:I 
*.PININFO en_samp_n:I en_samp_p:I en_update:I seq_comp:I seq_init:I seq_samp:I 
*.PININFO seq_update:I comp_out:O vdd_a:B vdd_d:B vdd_dac:B vin_n:B vin_p:B 
*.PININFO vss_a:B vss_d:B vss_dac:B
XXcapdriver_p_main dac_drive_botplate_main_p[15] dac_drive_botplate_main_p[14] 
+ dac_drive_botplate_main_p[13] dac_drive_botplate_main_p[12] 
+ dac_drive_botplate_main_p[11] dac_drive_botplate_main_p[10] 
+ dac_drive_botplate_main_p[9] dac_drive_botplate_main_p[8] 
+ dac_drive_botplate_main_p[7] dac_drive_botplate_main_p[6] 
+ dac_drive_botplate_main_p[5] dac_drive_botplate_main_p[4] 
+ dac_drive_botplate_main_p[3] dac_drive_botplate_main_p[2] 
+ dac_drive_botplate_main_p[1] dac_drive_botplate_main_p[0] dac_invert_p_main 
+ dac_state_p_main[15] dac_state_p_main[14] dac_state_p_main[13] 
+ dac_state_p_main[12] dac_state_p_main[11] dac_state_p_main[10] 
+ dac_state_p_main[9] dac_state_p_main[8] dac_state_p_main[7] 
+ dac_state_p_main[6] dac_state_p_main[5] dac_state_p_main[4] 
+ dac_state_p_main[3] dac_state_p_main[2] dac_state_p_main[1] 
+ dac_state_p_main[0] vdd_dac vss_dac / capdriver
XXcapdriver_p_diff dac_drive_botplate_diff_p[15] dac_drive_botplate_diff_p[14] 
+ dac_drive_botplate_diff_p[13] dac_drive_botplate_diff_p[12] 
+ dac_drive_botplate_diff_p[11] dac_drive_botplate_diff_p[10] 
+ dac_drive_botplate_diff_p[9] dac_drive_botplate_diff_p[8] 
+ dac_drive_botplate_diff_p[7] dac_drive_botplate_diff_p[6] 
+ dac_drive_botplate_diff_p[5] dac_drive_botplate_diff_p[4] 
+ dac_drive_botplate_diff_p[3] dac_drive_botplate_diff_p[2] 
+ dac_drive_botplate_diff_p[1] dac_drive_botplate_diff_p[0] dac_invert_p_diff 
+ dac_state_p_diff[15] dac_state_p_diff[14] dac_state_p_diff[13] 
+ dac_state_p_diff[12] dac_state_p_diff[11] dac_state_p_diff[10] 
+ dac_state_p_diff[9] dac_state_p_diff[8] dac_state_p_diff[7] 
+ dac_state_p_diff[6] dac_state_p_diff[5] dac_state_p_diff[4] 
+ dac_state_p_diff[3] dac_state_p_diff[2] dac_state_p_diff[1] 
+ dac_state_p_diff[0] vdd_dac vss_dac / capdriver
XXcapdriver_n_main dac_drive_botplate_main_n[15] dac_drive_botplate_main_n[14] 
+ dac_drive_botplate_main_n[13] dac_drive_botplate_main_n[12] 
+ dac_drive_botplate_main_n[11] dac_drive_botplate_main_n[10] 
+ dac_drive_botplate_main_n[9] dac_drive_botplate_main_n[8] 
+ dac_drive_botplate_main_n[7] dac_drive_botplate_main_n[6] 
+ dac_drive_botplate_main_n[5] dac_drive_botplate_main_n[4] 
+ dac_drive_botplate_main_n[3] dac_drive_botplate_main_n[2] 
+ dac_drive_botplate_main_n[1] dac_drive_botplate_main_n[0] dac_invert_n_main 
+ dac_state_n_main[15] dac_state_n_main[14] dac_state_n_main[13] 
+ dac_state_n_main[12] dac_state_n_main[11] dac_state_n_main[10] 
+ dac_state_n_main[9] dac_state_n_main[8] dac_state_n_main[7] 
+ dac_state_n_main[6] dac_state_n_main[5] dac_state_n_main[4] 
+ dac_state_n_main[3] dac_state_n_main[2] dac_state_n_main[1] 
+ dac_state_n_main[0] vdd_dac vss_dac / capdriver
XXcapdriver_n_diff dac_drive_botplate_diff_n[15] dac_drive_botplate_diff_n[14] 
+ dac_drive_botplate_diff_n[13] dac_drive_botplate_diff_n[12] 
+ dac_drive_botplate_diff_n[11] dac_drive_botplate_diff_n[10] 
+ dac_drive_botplate_diff_n[9] dac_drive_botplate_diff_n[8] 
+ dac_drive_botplate_diff_n[7] dac_drive_botplate_diff_n[6] 
+ dac_drive_botplate_diff_n[5] dac_drive_botplate_diff_n[4] 
+ dac_drive_botplate_diff_n[3] dac_drive_botplate_diff_n[2] 
+ dac_drive_botplate_diff_n[1] dac_drive_botplate_diff_n[0] dac_invert_n_diff 
+ dac_state_n_diff[15] dac_state_n_diff[14] dac_state_n_diff[13] 
+ dac_state_n_diff[12] dac_state_n_diff[11] dac_state_n_diff[10] 
+ dac_state_n_diff[9] dac_state_n_diff[8] dac_state_n_diff[7] 
+ dac_state_n_diff[6] dac_state_n_diff[5] dac_state_n_diff[4] 
+ dac_state_n_diff[3] dac_state_n_diff[2] dac_state_n_diff[1] 
+ dac_state_n_diff[0] vdd_dac vss_dac / capdriver
XXcaparray_p dac_drive_botplate_diff_p[15] dac_drive_botplate_diff_p[14] 
+ dac_drive_botplate_diff_p[13] dac_drive_botplate_diff_p[12] 
+ dac_drive_botplate_diff_p[11] dac_drive_botplate_diff_p[10] 
+ dac_drive_botplate_diff_p[9] dac_drive_botplate_diff_p[8] 
+ dac_drive_botplate_diff_p[7] dac_drive_botplate_diff_p[6] 
+ dac_drive_botplate_diff_p[5] dac_drive_botplate_diff_p[4] 
+ dac_drive_botplate_diff_p[3] dac_drive_botplate_diff_p[2] 
+ dac_drive_botplate_diff_p[1] dac_drive_botplate_diff_p[0] 
+ dac_drive_botplate_main_p[15] dac_drive_botplate_main_p[14] 
+ dac_drive_botplate_main_p[13] dac_drive_botplate_main_p[12] 
+ dac_drive_botplate_main_p[11] dac_drive_botplate_main_p[10] 
+ dac_drive_botplate_main_p[9] dac_drive_botplate_main_p[8] 
+ dac_drive_botplate_main_p[7] dac_drive_botplate_main_p[6] 
+ dac_drive_botplate_main_p[5] dac_drive_botplate_main_p[4] 
+ dac_drive_botplate_main_p[3] dac_drive_botplate_main_p[2] 
+ dac_drive_botplate_main_p[1] dac_drive_botplate_main_p[0] vss_a vdac_p / 
+ caparray
XXcaparray_n dac_drive_botplate_diff_n[15] dac_drive_botplate_diff_n[14] 
+ dac_drive_botplate_diff_n[13] dac_drive_botplate_diff_n[12] 
+ dac_drive_botplate_diff_n[11] dac_drive_botplate_diff_n[10] 
+ dac_drive_botplate_diff_n[9] dac_drive_botplate_diff_n[8] 
+ dac_drive_botplate_diff_n[7] dac_drive_botplate_diff_n[6] 
+ dac_drive_botplate_diff_n[5] dac_drive_botplate_diff_n[4] 
+ dac_drive_botplate_diff_n[3] dac_drive_botplate_diff_n[2] 
+ dac_drive_botplate_diff_n[1] dac_drive_botplate_diff_n[0] 
+ dac_drive_botplate_main_n[15] dac_drive_botplate_main_n[14] 
+ dac_drive_botplate_main_n[13] dac_drive_botplate_main_n[12] 
+ dac_drive_botplate_main_n[11] dac_drive_botplate_main_n[10] 
+ dac_drive_botplate_main_n[9] dac_drive_botplate_main_n[8] 
+ dac_drive_botplate_main_n[7] dac_drive_botplate_main_n[6] 
+ dac_drive_botplate_main_n[5] dac_drive_botplate_main_n[4] 
+ dac_drive_botplate_main_n[3] dac_drive_botplate_main_n[2] 
+ dac_drive_botplate_main_n[1] dac_drive_botplate_main_n[0] vss_a vdac_n / 
+ caparray
XXsampswitch_p clk_samp_p clk_samp_p_b vdd_a vin_p vdac_p vss_a / sampswitch
XXsampswitch_n clk_samp_n clk_samp_n_b vdd_a vin_n vdac_n vss_a / sampswitch
XXcomp clk_comp comp_out_n comp_out_p vdd_a vdac_n vdac_p vss_a / comp
XXadc_digital clk_comp clk_samp_n clk_samp_n_b clk_samp_p clk_samp_p_b 
+ comp_out comp_out_n comp_out_p dac_astate_n[15] dac_astate_n[14] 
+ dac_astate_n[13] dac_astate_n[12] dac_astate_n[11] dac_astate_n[10] 
+ dac_astate_n[9] dac_astate_n[8] dac_astate_n[7] dac_astate_n[6] 
+ dac_astate_n[5] dac_astate_n[4] dac_astate_n[3] dac_astate_n[2] 
+ dac_astate_n[1] dac_astate_n[0] dac_astate_p[15] dac_astate_p[14] 
+ dac_astate_p[13] dac_astate_p[12] dac_astate_p[11] dac_astate_p[10] 
+ dac_astate_p[9] dac_astate_p[8] dac_astate_p[7] dac_astate_p[6] 
+ dac_astate_p[5] dac_astate_p[4] dac_astate_p[3] dac_astate_p[2] 
+ dac_astate_p[1] dac_astate_p[0] dac_bstate_n[15] dac_bstate_n[14] 
+ dac_bstate_n[13] dac_bstate_n[12] dac_bstate_n[11] dac_bstate_n[10] 
+ dac_bstate_n[9] dac_bstate_n[8] dac_bstate_n[7] dac_bstate_n[6] 
+ dac_bstate_n[5] dac_bstate_n[4] dac_bstate_n[3] dac_bstate_n[2] 
+ dac_bstate_n[1] dac_bstate_n[0] dac_bstate_p[15] dac_bstate_p[14] 
+ dac_bstate_p[13] dac_bstate_p[12] dac_bstate_p[11] dac_bstate_p[10] 
+ dac_bstate_p[9] dac_bstate_p[8] dac_bstate_p[7] dac_bstate_p[6] 
+ dac_bstate_p[5] dac_bstate_p[4] dac_bstate_p[3] dac_bstate_p[2] 
+ dac_bstate_p[1] dac_bstate_p[0] dac_diffcaps dac_invert_n_diff 
+ dac_invert_n_main dac_invert_p_diff dac_invert_p_main dac_mode 
+ dac_state_n_diff[15] dac_state_n_diff[14] dac_state_n_diff[13] 
+ dac_state_n_diff[12] dac_state_n_diff[11] dac_state_n_diff[10] 
+ dac_state_n_diff[9] dac_state_n_diff[8] dac_state_n_diff[7] 
+ dac_state_n_diff[6] dac_state_n_diff[5] dac_state_n_diff[4] 
+ dac_state_n_diff[3] dac_state_n_diff[2] dac_state_n_diff[1] 
+ dac_state_n_diff[0] dac_state_n_main[15] dac_state_n_main[14] 
+ dac_state_n_main[13] dac_state_n_main[12] dac_state_n_main[11] 
+ dac_state_n_main[10] dac_state_n_main[9] dac_state_n_main[8] 
+ dac_state_n_main[7] dac_state_n_main[6] dac_state_n_main[5] 
+ dac_state_n_main[4] dac_state_n_main[3] dac_state_n_main[2] 
+ dac_state_n_main[1] dac_state_n_main[0] dac_state_p_diff[15] 
+ dac_state_p_diff[14] dac_state_p_diff[13] dac_state_p_diff[12] 
+ dac_state_p_diff[11] dac_state_p_diff[10] dac_state_p_diff[9] 
+ dac_state_p_diff[8] dac_state_p_diff[7] dac_state_p_diff[6] 
+ dac_state_p_diff[5] dac_state_p_diff[4] dac_state_p_diff[3] 
+ dac_state_p_diff[2] dac_state_p_diff[1] dac_state_p_diff[0] 
+ dac_state_p_main[15] dac_state_p_main[14] dac_state_p_main[13] 
+ dac_state_p_main[12] dac_state_p_main[11] dac_state_p_main[10] 
+ dac_state_p_main[9] dac_state_p_main[8] dac_state_p_main[7] 
+ dac_state_p_main[6] dac_state_p_main[5] dac_state_p_main[4] 
+ dac_state_p_main[3] dac_state_p_main[2] dac_state_p_main[1] 
+ dac_state_p_main[0] en_comp en_init en_samp_n en_samp_p en_update seq_comp 
+ seq_init seq_samp seq_update vdd_d vss_d / adc_digital
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    INVD3LVT
* View Name:    schematic
************************************************************************

.SUBCKT INVD3LVT I VDD VSS ZN
*.PININFO I:I ZN:O VDD:B VSS:B
MMU1_0-M_u2 ZN I VSS VSS nch_lvt l=60n w=390.0n m=1
MMU1_1-M_u2 ZN I VSS VSS nch_lvt l=60n w=390.0n m=1
MMU1_2-M_u2 ZN I VSS VSS nch_lvt l=60n w=390.0n m=1
MMU1_0-M_u3 ZN I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU1_1-M_u3 ZN I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU1_2-M_u3 ZN I VDD VDD pch_lvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    IND2D1LVT
* View Name:    schematic
************************************************************************

.SUBCKT IND2D1LVT A1 B1 VDD VSS ZN
*.PININFO A1:I B1:I ZN:O VDD:B VSS:B
MMI2-M_u3 net9 A1 VDD VDD pch_lvt l=60n w=260.0n m=1
MMI11 VDD B1 ZN VDD pch_lvt l=60n w=520.0n m=1
MM_u16 VDD net9 ZN VDD pch_lvt l=60n w=520.0n m=1
MMI13 net21 net9 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI2-M_u2 net9 A1 VSS VSS nch_lvt l=60n w=195.00n m=1
MMI12 ZN B1 net21 VSS nch_lvt l=60n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    CKND2LVT
* View Name:    schematic
************************************************************************

.SUBCKT CKND2LVT I VDD VSS ZN
*.PININFO I:I ZN:O VDD:B VSS:B
MM_u1_0 ZN I VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u1_1 ZN I VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2_1 ZN I VSS VSS nch_lvt l=60n w=310.0n m=1
MM_u2_0 ZN I VSS VSS nch_lvt l=60n w=310.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    ND3D1LVT
* View Name:    schematic
************************************************************************

.SUBCKT ND3D1LVT A1 A2 A3 VDD VSS ZN
*.PININFO A1:I A2:I A3:I ZN:O VDD:B VSS:B
MMI1-M_u5 net9 A2 net1 VSS nch_lvt l=60n w=390.0n m=1
MMI1-M_u4 ZN A1 net9 VSS nch_lvt l=60n w=390.0n m=1
MMI1-M_u6 net1 A3 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI1-M_u1 ZN A1 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI1-M_u3 ZN A3 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI1-M_u2 ZN A2 VDD VDD pch_lvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    ND2D1LVT
* View Name:    schematic
************************************************************************

.SUBCKT ND2D1LVT A1 A2 VDD VSS ZN
*.PININFO A1:I A2:I ZN:O VDD:B VSS:B
MMI1-M_u3 ZN A1 net1 VSS nch_lvt l=60n w=390.0n m=1
MMI1-M_u4 net1 A2 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI1-M_u1 ZN A1 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI1-M_u2 ZN A2 VDD VDD pch_lvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    NR2D2LVT
* View Name:    schematic
************************************************************************

.SUBCKT NR2D2LVT A1 A2 VDD VSS ZN
*.PININFO A1:I A2:I ZN:O VDD:B VSS:B
MMI1_1-M_u3 ZN A2 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI1_1-M_u4 ZN A1 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI1_0-M_u4 ZN A1 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI1_0-M_u3 ZN A2 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI1_1-M_u2 ZN A1 net17 VDD pch_lvt l=60n w=530.0n m=1
MMI1_0-M_u1 net25 A2 VDD VDD pch_lvt l=60n w=530.0n m=1
MMI1_0-M_u2 ZN A1 net25 VDD pch_lvt l=60n w=530.0n m=1
MMI1_1-M_u1 net17 A2 VDD VDD pch_lvt l=60n w=530.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    NR2XD1LVT
* View Name:    schematic
************************************************************************

.SUBCKT NR2XD1LVT A1 A2 VDD VSS ZN
*.PININFO A1:I A2:I ZN:O VDD:B VSS:B
MMI1-M_u3 ZN A2 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI1-M_u4 ZN A1 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI1-M_u1 net13 A2 VDD VDD pch_lvt l=60n w=1.04u m=1
MMI1-M_u2 ZN A1 net13 VDD pch_lvt l=60n w=1.04u m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    CKND2D1LVT
* View Name:    schematic
************************************************************************

.SUBCKT CKND2D1LVT A1 A2 VDD VSS ZN
*.PININFO A1:I A2:I ZN:O VDD:B VSS:B
MMI0-M_u3 ZN A1 net1 VSS nch_lvt l=60n w=390.0n m=1
MMI0-M_u4 net1 A2 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI0-M_u1 ZN A1 VDD VDD pch_lvt l=60n w=390.0n m=1
MMI0-M_u2 ZN A2 VDD VDD pch_lvt l=60n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    CKND2D2LVT
* View Name:    schematic
************************************************************************

.SUBCKT CKND2D2LVT A1 A2 VDD VSS ZN
*.PININFO A1:I A2:I ZN:O VDD:B VSS:B
MMI0_0-M_u1 ZN A1 VDD VDD pch_lvt l=60n w=390.0n m=1
MMI0_1-M_u2 ZN A2 VDD VDD pch_lvt l=60n w=390.0n m=1
MMI0_0-M_u2 ZN A2 VDD VDD pch_lvt l=60n w=390.0n m=1
MMI0_1-M_u1 ZN A1 VDD VDD pch_lvt l=60n w=390.0n m=1
MMI0_1-M_u4 net24 A2 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI0_0-M_u3 ZN A1 net17 VSS nch_lvt l=60n w=390.0n m=1
MMI0_1-M_u3 ZN A1 net24 VSS nch_lvt l=60n w=390.0n m=1
MMI0_0-M_u4 net17 A2 VSS VSS nch_lvt l=60n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    ND3D2LVT
* View Name:    schematic
************************************************************************

.SUBCKT ND3D2LVT A1 A2 A3 VDD VSS ZN
*.PININFO A1:I A2:I A3:I ZN:O VDD:B VSS:B
MMI0_0-M_u3 ZN A3 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI0_0-M_u1 ZN A1 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI0_1-M_u2 ZN A2 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI0_1-M_u3 ZN A3 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI0_0-M_u2 ZN A2 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI0_1-M_u1 ZN A1 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI0_1-M_u5 net44 A2 net37 VSS nch_lvt l=60n w=390.0n m=1
MMI0_1-M_u4 ZN A1 net44 VSS nch_lvt l=60n w=390.0n m=1
MMI0_1-M_u6 net37 A3 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI0_0-M_u6 net33 A3 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI0_0-M_u5 net29 A2 net33 VSS nch_lvt l=60n w=390.0n m=1
MMI0_0-M_u4 ZN A1 net29 VSS nch_lvt l=60n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    CKND1LVT
* View Name:    schematic
************************************************************************

.SUBCKT CKND1LVT I VDD VSS ZN
*.PININFO I:I ZN:O VDD:B VSS:B
MM_u2 ZN I VSS VSS nch_lvt l=60n w=310.0n m=1
MM_u1 ZN I VDD VDD pch_lvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    BUFFD16LVT
* View Name:    schematic
************************************************************************

.SUBCKT BUFFD16LVT I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
MMU8_0-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_3-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_9-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_5-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_6-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u2_3-M_u2 net123 I VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u2_1-M_u2 net123 I VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_13-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_4-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_1-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_14-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_12-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u2_4-M_u2 net123 I VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u2_2-M_u2 net123 I VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_11-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u2_0-M_u2 net123 I VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_15-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_8-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_2-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_7-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_10-M_u2 Z net123 VSS VSS nch_lvt l=60n w=390.0n m=1
MMU8_6-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_9-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_7-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_0-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2_1-M_u3 net123 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_4-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2_3-M_u3 net123 I VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2_0-M_u3 net123 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_14-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_12-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_11-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_8-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2_2-M_u3 net123 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_13-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2_4-M_u3 net123 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_1-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_2-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_3-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_5-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_10-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU8_15-M_u3 Z net123 VDD VDD pch_lvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    EDFCND2LVT
* View Name:    schematic
************************************************************************

.SUBCKT EDFCND2LVT CDN CP D E Q QN VDD VSS
*.PININFO CDN:I CP:I D:I E:I Q:O QN:O VDD:B VSS:B
MMI144-M_u1 net67 net20 VDD VDD pch_lvt l=60n w=400n m=1
MMI145-M_u3 Q net67 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI43 net81 net25 VDD VDD pch_lvt l=60n w=155.00n m=1
MMI149 net5 net79 net80 VDD pch_lvt l=60n w=340.0n m=1
MMI31-M_u3 net123 CP VDD VDD pch_lvt l=60n w=260.0n m=1
MMI29-M_u3 QN net161 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI27-M_u3 Q net67 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI146-M_u3 QN net161 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI147-M_u2 net67 CDN VDD VDD pch_lvt l=60n w=520.0n m=1
MMI44 net81 CDN VDD VDD pch_lvt l=60n w=150.0n m=1
MMI147-M_u1 net67 net20 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI17 net161 net125 net20 VDD pch_lvt l=60n w=150.0n m=1
MMI139 net80 D VDD VDD pch_lvt l=60n w=340.0n m=1
MMI138 net9 net125 net5 VDD pch_lvt l=60n w=340.0n m=1
MMI140 net33 net161 VDD VDD pch_lvt l=60n w=380.0n m=1
MMI151-M_u3 net161 net67 VDD VDD pch_lvt l=60n w=400n m=1
MMI13-M_u3 net25 net9 VDD VDD pch_lvt l=60n w=210.0n m=1
MMI150-M_u3 net125 net123 VDD VDD pch_lvt l=60n w=260.0n m=1
MMI16 net25 net123 net20 VDD pch_lvt l=60n w=390.0n m=1
MMI144-M_u2 net67 CDN VDD VDD pch_lvt l=60n w=400n m=1
MMI45 net9 net123 net81 VDD pch_lvt l=60n w=155.00n m=1
MMI141 net5 E net33 VDD pch_lvt l=60n w=380.0n m=1
MMI137-M_u3 net79 E VDD VDD pch_lvt l=60n w=290.0n m=1
MMI151-M_u2 net161 net67 VSS VSS nch_lvt l=60n w=270.0n m=1
MMI29-M_u2 QN net161 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI146-M_u2 QN net161 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI144-M_u4 net169 CDN VSS VSS nch_lvt l=60n w=200n m=1
MMI136 net124 net79 net149 VSS nch_lvt l=60n w=350.0n m=1
MMI18 net161 net123 net20 VSS nch_lvt l=60n w=150.0n m=1
MMI144-M_u3 net67 net20 net169 VSS nch_lvt l=60n w=200n m=1
MMI147-M_u3 net67 net20 net156 VSS nch_lvt l=60n w=200n m=1
MMI133 net149 net161 VSS VSS nch_lvt l=60n w=350.0n m=1
MMI145-M_u2 Q net67 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI137-M_u2 net79 E VSS VSS nch_lvt l=60n w=195.00n m=1
MMI13-M_u2 net25 net9 VSS VSS nch_lvt l=60n w=180.0n m=1
MMI135 net80 D VSS VSS nch_lvt l=60n w=210.0n m=1
MMI15 net25 net125 net20 VSS nch_lvt l=60n w=235.00n m=1
MMI150-M_u2 net125 net123 VSS VSS nch_lvt l=60n w=195.00n m=1
MMI132 net9 net123 net124 VSS nch_lvt l=60n w=290.0n m=1
MMI148 net124 E net80 VSS nch_lvt l=60n w=210.0n m=1
MMI31-M_u2 net123 CP VSS VSS nch_lvt l=60n w=195.00n m=1
MMI49 net104 CDN VSS VSS nch_lvt l=60n w=150.0n m=1
MMI147-M_u4 net156 CDN VSS VSS nch_lvt l=60n w=200n m=1
MMI48 net96 net25 net104 VSS nch_lvt l=60n w=150.0n m=1
MMI27-M_u2 Q net67 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI47 net9 net125 net96 VSS nch_lvt l=60n w=150.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    EDFCND4LVT
* View Name:    schematic
************************************************************************

.SUBCKT EDFCND4LVT CDN CP D E Q QN VDD VSS
*.PININFO CDN:I CP:I D:I E:I Q:O QN:O VDD:B VSS:B
MMI29-M_u2 QN net79 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI156-M_u2 net203 CP VSS VSS nch_lvt l=60n w=390.0n m=1
MMI144-M_u4 net97 CDN VSS VSS nch_lvt l=60n w=200n m=1
MMI136 net44 net95 net77 VSS nch_lvt l=60n w=350.0n m=1
MMI18 net79 net203 net83 VSS nch_lvt l=60n w=150.0n m=1
MMI151-M_u4 net64 CDN VSS VSS nch_lvt l=60n w=200n m=1
MMI144-M_u3 net11 net83 net97 VSS nch_lvt l=60n w=200n m=1
MMI133 net77 net79 VSS VSS nch_lvt l=60n w=350.0n m=1
MMI147-M_u2 QN net79 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI137-M_u2 net95 E VSS VSS nch_lvt l=60n w=195.00n m=1
MMI13-M_u2 net137 net5 VSS VSS nch_lvt l=60n w=190.0n m=1
MMI151-M_u3 net11 net83 net64 VSS nch_lvt l=60n w=200n m=1
MMI135 net32 D VSS VSS nch_lvt l=60n w=210.0n m=1
MMI15 net137 net33 net83 VSS nch_lvt l=60n w=235.00n m=1
MMI150-M_u2 Q net11 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI14-M_u2 net79 net11 VSS VSS nch_lvt l=60n w=465.00n m=1
MMI132 net5 net203 net44 VSS nch_lvt l=60n w=290.0n m=1
MMI155-M_u2 QN net79 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI32-M_u2 net33 net203 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI153 net44 E net32 VSS nch_lvt l=60n w=210.0n m=1
MMI149-M_u2 Q net11 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI49 net21 CDN VSS VSS nch_lvt l=60n w=150.0n m=1
MMI48 net8 net137 net21 VSS nch_lvt l=60n w=150.0n m=1
MMI27-M_u2 Q net11 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI154-M_u2 Q net11 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI47 net5 net33 net8 VSS nch_lvt l=60n w=150.0n m=1
MMI148-M_u2 QN net79 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI151-M_u2 net11 CDN VDD VDD pch_lvt l=60n w=520.0n m=1
MMI14-M_u3 net79 net11 VDD VDD pch_lvt l=60n w=660.0n m=1
MMI144-M_u1 net11 net83 VDD VDD pch_lvt l=60n w=400n m=1
MMI32-M_u3 net33 net203 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI43 net128 net137 VDD VDD pch_lvt l=60n w=155.00n m=1
MMI29-M_u3 QN net79 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI27-M_u3 Q net11 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI147-M_u3 QN net79 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI44 net128 CDN VDD VDD pch_lvt l=60n w=150.0n m=1
MMI17 net79 net33 net83 VDD pch_lvt l=60n w=150.0n m=1
MMI139 net32 D VDD VDD pch_lvt l=60n w=340.0n m=1
MMI138 net5 net33 net141 VDD pch_lvt l=60n w=340.0n m=1
MMI151-M_u1 net11 net83 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI140 net124 net79 VDD VDD pch_lvt l=60n w=380.0n m=1
MMI156-M_u3 net203 CP VDD VDD pch_lvt l=60n w=520.0n m=1
MMI13-M_u3 net137 net5 VDD VDD pch_lvt l=60n w=210.0n m=1
MMI150-M_u3 Q net11 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI149-M_u3 Q net11 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI152 net141 net95 net32 VDD pch_lvt l=60n w=340.0n m=1
MMI16 net137 net203 net83 VDD pch_lvt l=60n w=390.0n m=1
MMI154-M_u3 Q net11 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI144-M_u2 net11 CDN VDD VDD pch_lvt l=60n w=400n m=1
MMI45 net5 net203 net128 VDD pch_lvt l=60n w=155.00n m=1
MMI141 net141 E net124 VDD pch_lvt l=60n w=380.0n m=1
MMI137-M_u3 net95 E VDD VDD pch_lvt l=60n w=260.0n m=1
MMI148-M_u3 QN net79 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI155-M_u3 QN net79 VDD VDD pch_lvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    BUFFD6LVT
* View Name:    schematic
************************************************************************

.SUBCKT BUFFD6LVT I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
MM_u3_1-M_u2 Z net9 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u3_2-M_u2 Z net9 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u3_3-M_u2 Z net9 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u2_1-M_u2 net9 I VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u3_0-M_u2 Z net9 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u2_0-M_u2 net9 I VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u3_4-M_u2 Z net9 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u3_5-M_u2 Z net9 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u3_4-M_u3 Z net9 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_0-M_u3 Z net9 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_5-M_u3 Z net9 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2_1-M_u3 net9 I VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2_0-M_u3 net9 I VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_2-M_u3 Z net9 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_1-M_u3 Z net9 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_3-M_u3 Z net9 VDD VDD pch_lvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    CKBD16LVT
* View Name:    schematic
************************************************************************

.SUBCKT CKBD16LVT I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
DDI3 VSS I ndio_lvt area=6.6e-14 pj=1.18e-06 m=1
MMU21_12 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_4 net5 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_15 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_7 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_0 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_1 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_11 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_5 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_3 net5 I VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_0 net5 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_10 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_13 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_3 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_4 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_2 net5 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_6 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_9 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_8 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_1 net5 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_2 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_14 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU23_7 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MM_u15_3 net5 I VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_5 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_10 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_12 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_4 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MM_u15_4 net5 I VSS VSS nch_lvt l=60n w=310.0n m=1
MM_u15_1 net5 I VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_15 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_1 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_8 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_6 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_13 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_11 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MM_u15_2 net5 I VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_9 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_3 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_0 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_14 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_2 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MM_u15_0 net5 I VSS VSS nch_lvt l=60n w=310.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    CKBD3LVT
* View Name:    schematic
************************************************************************

.SUBCKT CKBD3LVT I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
MMU23_1 Z net9 VSS VSS nch_lvt l=60n w=310.0n m=1
MM_u15 net9 I VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_0 Z net9 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_2 Z net9 VSS VSS nch_lvt l=60n w=310.0n m=1
MM_u3 net9 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_0 Z net9 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_1 Z net9 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_2 Z net9 VDD VDD pch_lvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    BUFFD3LVT
* View Name:    schematic
************************************************************************

.SUBCKT BUFFD3LVT I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
MM_u3_0-M_u3 Z net11 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_2-M_u3 Z net11 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_1-M_u3 Z net11 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2-M_u3 net11 I VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_1-M_u2 Z net11 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u3_2-M_u2 Z net11 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u2-M_u2 net11 I VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u3_0-M_u2 Z net11 VSS VSS nch_lvt l=60n w=390.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    CKBD4LVT
* View Name:    schematic
************************************************************************

.SUBCKT CKBD4LVT I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
MM_u15_1 net11 I VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_1 Z net11 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_3 Z net11 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_0 Z net11 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_2 Z net11 VSS VSS nch_lvt l=60n w=310.0n m=1
MM_u15_0 net11 I VSS VSS nch_lvt l=60n w=310.0n m=1
MMU21_0 Z net11 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_1 Z net11 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_0 net11 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_3 Z net11 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_1 net11 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_2 Z net11 VDD VDD pch_lvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    CKBD8LVT
* View Name:    schematic
************************************************************************

.SUBCKT CKBD8LVT I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
DDI3 VSS I ndio_lvt area=6.6e-14 pj=1.18e-06 m=1
MMU21_7 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_0 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_1 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_5 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_0 net5 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_3 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_4 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_2 net5 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_6 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_1 net5 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_2 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU23_7 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_5 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_4 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_1 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MM_u15 net5 I VSS VSS nch_lvt l=60n w=780.0n m=1
MMU23_6 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_3 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_0 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_2 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    DEL4LVT
* View Name:    schematic
************************************************************************

.SUBCKT DEL4LVT I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
MMI4-M_u3 net11 net13 VDD VDD pch_lvt l=1u w=300n m=1
MMI7-M_u3 net25 net9 VDD VDD pch_lvt l=1u w=300n m=1
MMI5-M_u3 net13 net47 VDD VDD pch_lvt l=1u w=300n m=1
MMI8-M_u3 net9 net11 VDD VDD pch_lvt l=1u w=300n m=1
MMI3-M_u3 Z net25 VDD VDD pch_lvt l=60n w=520.0n m=1
MMI6-M_u3 net47 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMI5-M_u2 net13 net47 VSS VSS nch_lvt l=1u w=300n m=1
MMI8-M_u2 net9 net11 VSS VSS nch_lvt l=1u w=300n m=1
MMI3-M_u2 Z net25 VSS VSS nch_lvt l=60n w=390.0n m=1
MMI4-M_u2 net11 net13 VSS VSS nch_lvt l=1u w=300n m=1
MMI6-M_u2 net47 I VSS VSS nch_lvt l=60n w=390.0n m=1
MMI7-M_u2 net25 net9 VSS VSS nch_lvt l=1u w=300n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    CKBD1LVT
* View Name:    schematic
************************************************************************

.SUBCKT CKBD1LVT I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
MM_u15 net5 I VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MM_u3 net5 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    BUFFD8LVT
* View Name:    schematic
************************************************************************

.SUBCKT BUFFD8LVT I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
MM_u7_5-M_u2 Z net67 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u7_1-M_u2 Z net67 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u7_0-M_u2 Z net67 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u2_1-M_u2 net67 I VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u7_6-M_u2 Z net67 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u7_3-M_u2 Z net67 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u2_2-M_u2 net67 I VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u2_0-M_u2 net67 I VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u7_2-M_u2 Z net67 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u7_7-M_u2 Z net67 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u7_4-M_u2 Z net67 VSS VSS nch_lvt l=60n w=390.0n m=1
MM_u7_0-M_u3 Z net67 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u7_4-M_u3 Z net67 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u7_3-M_u3 Z net67 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2_1-M_u3 net67 I VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u7_5-M_u3 Z net67 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u7_1-M_u3 Z net67 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2_0-M_u3 net67 I VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u2_2-M_u3 net67 I VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u7_6-M_u3 Z net67 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u7_2-M_u3 Z net67 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u7_7-M_u3 Z net67 VDD VDD pch_lvt l=60n w=520.0n m=1
.ENDS

************************************************************************
* Library Name: tcbn65lplvt
* Cell Name:    CKBD6LVT
* View Name:    schematic
************************************************************************

.SUBCKT CKBD6LVT I VDD VSS Z
*.PININFO I:I Z:O VDD:B VSS:B
DDI3 VSS I ndio_lvt area=6.6e-14 pj=1.18e-06 m=1
MMU21_0 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_1 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_5 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_0 net5 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_3 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_4 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MM_u3_1 net5 I VDD VDD pch_lvt l=60n w=520.0n m=1
MMU21_2 Z net5 VDD VDD pch_lvt l=60n w=520.0n m=1
MMU23_5 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_4 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_1 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MM_u15 net5 I VSS VSS nch_lvt l=60n w=520.0n m=1
MMU23_3 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_0 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
MMU23_2 Z net5 VSS VSS nch_lvt l=60n w=310.0n m=1
.ENDS

************************************************************************
* Library Name: frida
* Cell Name:    frida_core
* View Name:    schematic
************************************************************************

.SUBCKT frida_core comp_out reset_b seq_comp seq_init seq_logic seq_samp 
+ spi_cs_b spi_sclk spi_sdi spi_sdo vdd_a vdd_d vdd_dac vin_n vin_p vss_a 
+ vss_d vss_dac
*.PININFO reset_b:I seq_comp:I seq_init:I seq_logic:I seq_samp:I spi_cs_b:I 
*.PININFO spi_sclk:I spi_sdi:I vin_n:I vin_p:I comp_out:O spi_sdo:O vdd_a:B 
*.PININFO vdd_d:B vdd_dac:B vss_a:B vss_d:B vss_dac:B
XXadc_array_adc_inst[10] adc_comparator_out[10] net2549 net2550 net2554 
+ net2556 net2557 net2559 net2561 net2563 net2564 net2566 net2569 net2571 
+ net2573 net2575 net2577 net2588 net2488 net2490 net2491 net2494 net2497 
+ net2499 net2501 net2503 net2505 net2506 net2508 net2511 net2513 net2515 
+ net2520 net2522 net2589 net2591 net2608 net2619 net2633 net2646 net2469 
+ net2481 net2483 net2485 net2495 net2517 net2537 net2553 net2572 net2657 
+ net2523 net2524 net2526 net2529 net2531 net2532 net2533 net2535 net2539 
+ net2541 net2542 net2543 net2544 net2546 net2547 net2548 net2607 net2609 
+ net2611 net2614 net2612 net2613 net2610 net2846 net2816 net2832 net2862 
+ vdd_a vdd_d vdd_dac vin_n vin_p vss_a vss_d vss_dac / adc
XXadc_array_adc_inst[11] adc_comparator_out[11] net2549 net2550 net2554 
+ net2556 net2557 net2559 net2561 net2563 net2564 net2566 net2569 net2571 
+ net2573 net2575 net2577 net2588 net2488 net2490 net2491 net2494 net2497 
+ net2499 net2501 net2503 net2505 net2506 net2508 net2511 net2513 net2515 
+ net2520 net2522 net2589 net2591 net2608 net2619 net2633 net2646 net2469 
+ net2481 net2483 net2485 net2495 net2518 net2538 net2553 net2572 net2657 
+ net2523 net2524 net2526 net2529 net2531 net2532 net2533 net2535 net2539 
+ net2541 net2542 net2543 net2544 net2546 net2547 net2548 net2600 net2601 
+ net2603 net2606 net2604 net2605 net2602 net2845 net2815 net2831 net2861 
+ vdd_a vdd_d vdd_dac vin_n vin_p vss_a vss_d vss_dac / adc
XXadc_array_adc_inst[4] adc_comparator_out[4] net2549 net2551 net2555 net2556 
+ net2557 net2558 net2560 net2562 net2565 net2567 net2568 net2570 net2574 
+ net2576 net2578 net2587 net2489 net2490 net2492 net2493 net2496 net2498 
+ net2500 net2502 net2504 net2507 net2509 net2510 net2512 net2514 net2519 
+ net2521 net2589 net2591 net2608 net2619 net2632 net2646 net2469 net2481 
+ net2482 net2486 net2495 net2517 net2537 net2552 net2572 net2657 net2523 
+ net2525 net2527 net2528 net2530 net2532 net2533 net2534 net2539 net2540 
+ net2542 net2543 net2544 net2545 net2547 net2548 net2471 net2472 net2474 
+ net2478 net2475 net2476 net2473 net2843 net2813 net2829 net2859 vdd_a vdd_d 
+ vdd_dac vin_n vin_p vss_a vss_d vss_dac / adc
XXadc_array_adc_inst[7] adc_comparator_out[7] net2549 net2550 net2554 net2556 
+ net2557 net2559 net2561 net2563 net2564 net2566 net2569 net2571 net2573 
+ net2575 net2577 net2588 net2488 net2490 net2491 net2494 net2497 net2499 
+ net2501 net2503 net2505 net2506 net2508 net2511 net2513 net2515 net2520 
+ net2522 net2589 net2591 net2608 net2619 net2633 net2646 net2469 net2481 
+ net2483 net2485 net2495 net2518 net2538 net2553 net2572 net2657 net2523 
+ net2524 net2526 net2529 net2531 net2532 net2533 net2535 net2539 net2541 
+ net2542 net2543 net2544 net2546 net2547 net2548 net2636 net2637 net2639 
+ net2642 net2640 net2641 net2638 net2839 net2809 net2825 net2855 vdd_a vdd_d 
+ vdd_dac vin_n vin_p vss_a vss_d vss_dac / adc
XXadc_array_adc_inst[8] adc_comparator_out[8] net2549 net2551 net2555 net2556 
+ net2557 net2558 net2560 net2562 net2565 net2567 net2568 net2570 net2574 
+ net2576 net2578 net2587 net2489 net2490 net2492 net2493 net2496 net2498 
+ net2500 net2502 net2504 net2507 net2509 net2510 net2512 net2514 net2519 
+ net2521 net2589 net2591 net2608 net2619 net2632 net2646 net2469 net2481 
+ net2482 net2486 net2495 net2517 net2537 net2552 net2572 net2657 net2523 
+ net2525 net2527 net2528 net2530 net2532 net2533 net2534 net2539 net2540 
+ net2542 net2543 net2544 net2545 net2547 net2548 net2624 net2625 net2627 
+ net2631 net2628 net2629 net2626 net2848 net2818 net2834 net2864 vdd_a vdd_d 
+ vdd_dac vin_n vin_p vss_a vss_d vss_dac / adc
XXadc_array_adc_inst[5] adc_comparator_out[5] net2549 net2551 net2555 net2556 
+ net2557 net2558 net2560 net2562 net2565 net2567 net2568 net2570 net2574 
+ net2576 net2578 net2587 net2488 net2490 net2492 net2493 net2496 net2498 
+ net2500 net2502 net2504 net2507 net2509 net2510 net2512 net2514 net2519 
+ net2521 net2589 net2591 net2608 net2619 net2632 net2646 net2469 net2481 
+ net2482 net2486 net2495 net2517 net2537 net2552 net2572 net2657 net2523 
+ net2525 net2527 net2528 net2530 net2532 net2533 net2534 net2539 net2540 
+ net2542 net2543 net2544 net2545 net2547 net2548 net2651 net2652 net2654 
+ net2470 net2655 net2656 net2653 net2843 net2813 net2829 net2859 vdd_a vdd_d 
+ vdd_dac vin_n vin_p vss_a vss_d vss_dac / adc
XXadc_array_adc_inst[6] adc_comparator_out[6] net2549 net2550 net2554 net2556 
+ net2557 net2559 net2561 net2563 net2564 net2566 net2569 net2571 net2573 
+ net2575 net2577 net2588 net2488 net2490 net2491 net2494 net2497 net2499 
+ net2501 net2503 net2505 net2506 net2508 net2511 net2513 net2515 net2520 
+ net2522 net2589 net2591 net2608 net2619 net2633 net2646 net2469 net2481 
+ net2483 net2485 net2495 net2517 net2537 net2553 net2572 net2657 net2523 
+ net2524 net2526 net2529 net2531 net2532 net2533 net2535 net2539 net2541 
+ net2542 net2543 net2544 net2546 net2547 net2548 net2643 net2644 net2647 
+ net2650 net2648 net2649 net2645 net2840 net2810 net2826 net2856 vdd_a vdd_d 
+ vdd_dac vin_n vin_p vss_a vss_d vss_dac / adc
XXadc_array_adc_inst[9] adc_comparator_out[9] net2549 net2551 net2555 net2556 
+ net2557 net2558 net2560 net2562 net2565 net2567 net2568 net2570 net2574 
+ net2576 net2578 net2587 net2488 net2490 net2492 net2493 net2496 net2498 
+ net2500 net2502 net2504 net2507 net2509 net2510 net2512 net2514 net2519 
+ net2521 net2589 net2591 net2608 net2619 net2632 net2646 net2469 net2481 
+ net2482 net2486 net2495 net2517 net2537 net2552 net2572 net2657 net2523 
+ net2525 net2527 net2528 net2530 net2532 net2533 net2534 net2539 net2540 
+ net2542 net2543 net2544 net2545 net2547 net2548 net2615 net2616 net2618 
+ net2623 net2620 net2621 net2617 net2848 net2818 net2834 net2864 vdd_a vdd_d 
+ vdd_dac vin_n vin_p vss_a vss_d vss_dac / adc
XXadc_array_adc_inst[12] adc_comparator_out[12] net2549 net2551 net2555 
+ net2556 net2557 net2558 net2560 net2562 net2565 net2567 net2568 net2570 
+ net2574 net2576 net2578 net2587 net2489 net2490 net2492 net2493 net2496 
+ net2498 net2500 net2502 net2504 net2507 net2509 net2510 net2512 net2514 
+ net2519 net2521 net2589 net2591 net2608 net2619 net2632 net2646 net2469 
+ net2481 net2482 net2486 net2495 net2517 net2537 net2552 net2572 net2657 
+ net2523 net2525 net2527 net2528 net2530 net2532 net2533 net2534 net2539 
+ net2540 net2542 net2543 net2544 net2545 net2547 net2548 spi_bits[154] 
+ spi_bits[153] spi_bits[151] net2597 spi_bits[150] spi_bits[149] 
+ spi_bits[152] net2849 net2819 net2835 net2865 vdd_a vdd_d vdd_dac vin_n 
+ vin_p vss_a vss_d vss_dac / adc
XXadc_array_adc_inst[0] adc_comparator_out[0] net2549 net2551 net2555 net2556 
+ net2557 net2558 net2560 net2562 net2565 net2567 net2568 net2570 net2574 
+ net2576 net2578 net2587 net2489 net2490 net2492 net2493 net2496 net2498 
+ net2500 net2502 net2504 net2507 net2509 net2510 net2512 net2514 net2519 
+ net2521 net2589 net2591 net2608 net2619 net2632 net2646 net2469 net2481 
+ net2482 net2486 net2495 net2517 net2537 net2552 net2572 net2657 net2523 
+ net2525 net2527 net2528 net2530 net2532 net2533 net2534 net2539 net2540 
+ net2542 net2543 net2544 net2545 net2547 net2548 spi_bits[70] spi_bits[69] 
+ spi_bits[67] spi_bits[64] spi_bits[66] spi_bits[65] spi_bits[68] net2842 
+ net2812 net2828 net2858 vdd_a vdd_d vdd_dac vin_n vin_p vss_a vss_d vss_dac 
+ / adc
XXadc_array_adc_inst[13] adc_comparator_out[13] net2549 net2551 net2555 
+ net2556 net2557 net2558 net2560 net2562 net2565 net2567 net2568 net2570 
+ net2574 net2576 net2578 net2587 net2488 net2490 net2492 net2493 net2496 
+ net2498 net2500 net2502 net2504 net2507 net2509 net2510 net2512 net2514 
+ net2519 net2521 net2589 net2591 net2608 net2619 net2632 net2646 net2469 
+ net2481 net2482 net2486 net2495 net2517 net2537 net2552 net2572 net2657 
+ net2523 net2525 net2527 net2528 net2530 net2532 net2533 net2534 net2539 
+ net2540 net2542 net2543 net2544 net2545 net2547 net2548 spi_bits[161] 
+ spi_bits[160] spi_bits[158] net2590 spi_bits[157] spi_bits[156] 
+ spi_bits[159] net2849 net2819 net2835 net2865 vdd_a vdd_d vdd_dac vin_n 
+ vin_p vss_a vss_d vss_dac / adc
XXadc_array_adc_inst[14] adc_comparator_out[14] net2549 net2550 net2554 
+ net2556 net2557 net2559 net2561 net2563 net2564 net2566 net2569 net2571 
+ net2573 net2575 net2577 net2588 net2488 net2490 net2491 net2494 net2497 
+ net2499 net2501 net2503 net2505 net2506 net2508 net2511 net2513 net2515 
+ net2520 net2522 net2589 net2591 net2608 net2619 net2633 net2646 net2469 
+ net2481 net2483 net2485 net2495 net2517 net2537 net2553 net2572 net2657 
+ net2523 net2524 net2526 net2529 net2531 net2532 net2533 net2535 net2539 
+ net2541 net2542 net2543 net2544 net2546 net2547 net2548 spi_bits[168] 
+ spi_bits[167] spi_bits[165] spi_bits[162] spi_bits[164] spi_bits[163] 
+ spi_bits[166] net2847 net2817 net2833 net2863 vdd_a vdd_d vdd_dac vin_n 
+ vin_p vss_a vss_d vss_dac / adc
XXadc_array_adc_inst[15] adc_comparator_out[15] net2549 net2550 net2554 
+ net2556 net2557 net2559 net2561 net2563 net2564 net2566 net2569 net2571 
+ net2573 net2575 net2577 net2588 net2488 net2490 net2491 net2494 net2497 
+ net2499 net2501 net2503 net2505 net2506 net2508 net2511 net2513 net2515 
+ net2520 net2522 net2589 net2591 net2608 net2619 net2633 net2646 net2469 
+ net2481 net2483 net2485 net2495 net2518 net2538 net2553 net2572 net2657 
+ net2523 net2524 net2526 net2529 net2531 net2532 net2533 net2535 net2539 
+ net2541 net2542 net2543 net2544 net2546 net2547 net2548 spi_bits[175] 
+ spi_bits[174] spi_bits[172] spi_bits[169] spi_bits[171] spi_bits[170] 
+ spi_bits[173] net2845 net2815 net2831 net2861 vdd_a vdd_d vdd_dac vin_n 
+ vin_p vss_a vss_d vss_dac / adc
XXadc_array_adc_inst[1] adc_comparator_out[1] net2549 net2551 net2555 net2556 
+ net2557 net2558 net2560 net2562 net2565 net2567 net2568 net2570 net2574 
+ net2576 net2578 net2587 net2488 net2490 net2492 net2493 net2496 net2498 
+ net2500 net2502 net2504 net2507 net2509 net2510 net2512 net2514 net2519 
+ net2521 net2589 net2591 net2608 net2619 net2632 net2646 net2469 net2481 
+ net2482 net2486 net2495 net2517 net2537 net2552 net2572 net2660 net2523 
+ net2525 net2527 net2528 net2530 net2532 net2533 net2534 net2539 net2540 
+ net2542 net2543 net2544 net2545 net2547 net2548 spi_bits[77] spi_bits[76] 
+ spi_bits[74] net2484 spi_bits[73] spi_bits[72] spi_bits[75] net2842 net2812 
+ net2828 net2858 vdd_a vdd_d vdd_dac vin_n vin_p vss_a vss_d vss_dac / adc
XXadc_array_adc_inst[2] adc_comparator_out[2] net2549 net2550 net2554 net2556 
+ net2557 net2559 net2561 net2563 net2564 net2566 net2569 net2571 net2573 
+ net2575 net2577 net2588 net2488 net2490 net2491 net2494 net2497 net2499 
+ net2501 net2503 net2505 net2506 net2508 net2511 net2513 net2515 net2520 
+ net2522 net2589 net2591 net2608 net2619 net2633 net2646 net2469 net2481 
+ net2483 net2485 net2495 net2517 net2537 net2553 net2572 net2660 net2523 
+ net2524 net2526 net2529 net2531 net2532 net2533 net2535 net2539 net2541 
+ net2542 net2543 net2544 net2546 net2547 net2548 spi_bits[84] spi_bits[83] 
+ spi_bits[81] spi_bits[78] spi_bits[80] spi_bits[79] spi_bits[82] net2841 
+ net2811 net2827 net2857 vdd_a vdd_d vdd_dac vin_n vin_p vss_a vss_d vss_dac 
+ / adc
XXadc_array_adc_inst[3] adc_comparator_out[3] net2549 net2550 net2554 net2556 
+ net2557 net2559 net2561 net2563 net2564 net2566 net2569 net2571 net2573 
+ net2575 net2577 net2588 net2488 net2490 net2491 net2494 net2497 net2499 
+ net2501 net2503 net2505 net2506 net2508 net2511 net2513 net2515 net2520 
+ net2522 net2589 net2591 net2608 net2619 net2633 net2646 net2469 net2481 
+ net2483 net2485 net2495 net2518 net2538 net2553 net2572 net2660 net2523 
+ net2524 net2526 net2529 net2531 net2532 net2533 net2535 net2539 net2541 
+ net2542 net2543 net2544 net2546 net2547 net2548 spi_bits[91] spi_bits[90] 
+ spi_bits[88] spi_bits[85] spi_bits[87] spi_bits[86] spi_bits[89] net2839 
+ net2809 net2825 net2855 vdd_a vdd_d vdd_dac vin_n vin_p vss_a vss_d vss_dac 
+ / adc
XXcomp_mux_43_ net2580 vdd_d vss_d comp_mux_00_ / INVD3LVT
XXclkload4 clknet_4_9_leaf_spi_sclk vdd_d vss_d _unconnected_187 / INVD3LVT
XXcomp_mux_44_ net2756 net2468 vdd_d vss_d comp_mux_01_ / IND2D1LVT
XXcomp_mux_46_ net2752 net2581 vdd_d vss_d comp_mux_03_ / IND2D1LVT
XXcomp_mux_49_ net2749 comp_mux_00_ vdd_d vss_d comp_mux_06_ / IND2D1LVT
XXcomp_mux_60_ net2759 net2579 vdd_d vss_d comp_mux_17_ / IND2D1LVT
XXcomp_mux_65_ adc_comparator_out[1] net2581 vdd_d vss_d comp_mux_22_ / 
+ IND2D1LVT
XXcomp_mux_81_ net2734 net2580 vdd_d vss_d comp_mux_38_ / IND2D1LVT
XXinput1 reset_b vdd_d vss_d net1 / BUFFD2LVT
XXinput2 spi_cs_b vdd_d vss_d net2 / BUFFD2LVT
XXinput3 spi_sdi vdd_d vss_d net3 / BUFFD2LVT
XXoutput4 net4 vdd_d vss_d comp_out / BUFFD2LVT
XXplace2585 net2584 vdd_d vss_d net2585 / BUFFD2LVT
XXplace2634 spi_bits[119] vdd_d vss_d net2634 / BUFFD2LVT
XXplace2598 spi_bits[147] vdd_d vss_d net2598 / BUFFD2LVT
XXplace2697 net2696 vdd_d vss_d net2697 / BUFFD2LVT
XXplace2727 net2726 vdd_d vss_d net2727 / BUFFD2LVT
XXplace2731 net2730 vdd_d vss_d net2731 / BUFFD2LVT
XXplace2733 net2894 vdd_d vss_d net2733 / BUFFD2LVT
XXplace2666 net2665 vdd_d vss_d net2666 / BUFFD2LVT
XXplace2691 comp_mux_23_ vdd_d vss_d net2691 / BUFFD2LVT
XXplace2466 net5 vdd_d vss_d net2466 / BUFFD2LVT
XXplace2744 net2743 vdd_d vss_d net2744 / BUFFD2LVT
XXplace2740 net2739 vdd_d vss_d net2740 / BUFFD2LVT
XXplace2735 net2893 vdd_d vss_d net2735 / BUFFD2LVT
XXplace2737 net2892 vdd_d vss_d net2737 / BUFFD2LVT
XXplace2748 net2747 vdd_d vss_d net2748 / BUFFD2LVT
XXplace2751 net2750 vdd_d vss_d net2751 / BUFFD2LVT
XXplace2755 net2754 vdd_d vss_d net2755 / BUFFD2LVT
XXplace2758 net2757 vdd_d vss_d net2758 / BUFFD2LVT
XXplace2761 net2760 vdd_d vss_d net2761 / BUFFD2LVT
XXcomp_mux_47_ spi_bits[177] vdd_d vss_d comp_mux_04_ / CKND2LVT
XXcomp_mux_48_ comp_mux_01_ comp_mux_03_ comp_mux_04_ vdd_d vss_d comp_mux_05_ 
+ / ND3D1LVT
XXcomp_mux_52_ comp_mux_06_ comp_mux_08_ spi_bits[177] vdd_d vss_d 
+ comp_mux_09_ / ND3D1LVT
XXcomp_mux_53_ comp_mux_05_ comp_mux_09_ spi_bits[178] vdd_d vss_d 
+ comp_mux_10_ / ND3D1LVT
XXcomp_mux_63_ comp_mux_14_ comp_mux_18_ comp_mux_19_ vdd_d vss_d comp_mux_20_ 
+ / ND3D1LVT
XXcomp_mux_64_ comp_mux_10_ comp_mux_20_ spi_bits[179] vdd_d vss_d 
+ comp_mux_21_ / ND3D1LVT
XXcomp_mux_68_ comp_mux_22_ comp_mux_24_ comp_mux_04_ vdd_d vss_d comp_mux_25_ 
+ / ND3D1LVT
XXcomp_mux_73_ comp_mux_27_ comp_mux_29_ spi_bits[177] vdd_d vss_d 
+ comp_mux_30_ / ND3D1LVT
XXcomp_mux_74_ comp_mux_25_ comp_mux_30_ comp_mux_19_ vdd_d vss_d comp_mux_31_ 
+ / ND3D1LVT
XXcomp_mux_50_ net2745 vdd_d vss_d comp_mux_07_ / CKND0LVT
XXcomp_mux_62_ spi_bits[178] vdd_d vss_d comp_mux_19_ / CKND0LVT
XXcomp_mux_66_ adc_comparator_out[0] vdd_d vss_d comp_mux_23_ / CKND0LVT
XXcomp_mux_69_ adc_comparator_out[2] vdd_d vss_d comp_mux_26_ / CKND0LVT
XXcomp_mux_71_ adc_comparator_out[3] vdd_d vss_d comp_mux_28_ / CKND0LVT
XXcomp_mux_84_ spi_bits[179] vdd_d vss_d comp_mux_41_ / CKND0LVT
XXcomp_mux_51_ comp_mux_07_ net2881 vdd_d vss_d comp_mux_08_ / ND2D1LVT
XXcomp_mux_67_ net2691 net2468 vdd_d vss_d comp_mux_24_ / ND2D1LVT
XXcomp_mux_77_ comp_mux_32_ comp_mux_33_ vdd_d vss_d comp_mux_34_ / ND2D1LVT
XXcomp_mux_82_ comp_mux_37_ comp_mux_38_ vdd_d vss_d comp_mux_39_ / ND2D1LVT
XXcomp_mux_86_ comp_mux_21_ comp_mux_42_ vdd_d vss_d net4 / ND2D1LVT
XXcomp_mux_54_ net2468 net2732 vdd_d vss_d comp_mux_11_ / ND2D2LVT
XXcomp_mux_55_ net2581 net2728 vdd_d vss_d comp_mux_12_ / ND2D2LVT
XXcomp_mux_56_ comp_mux_11_ comp_mux_12_ vdd_d vss_d comp_mux_13_ / ND2D2LVT
XXcomp_mux_57_ comp_mux_13_ comp_mux_04_ vdd_d vss_d comp_mux_14_ / ND2D2LVT
XXcomp_mux_61_ comp_mux_16_ comp_mux_17_ vdd_d vss_d comp_mux_18_ / ND2D2LVT
XXcomp_mux_75_ net2468 net2741 vdd_d vss_d comp_mux_32_ / ND2D2LVT
XXcomp_mux_58_ net2580 net2762 vdd_d vss_d comp_mux_15_ / NR2D2LVT
XXcomp_mux_79_ net2580 net2736 vdd_d vss_d comp_mux_36_ / NR2D2LVT
XXcomp_mux_59_ comp_mux_15_ comp_mux_04_ vdd_d vss_d comp_mux_16_ / NR2XD1LVT
XXcomp_mux_80_ comp_mux_36_ comp_mux_04_ vdd_d vss_d comp_mux_37_ / NR2XD1LVT
XXcomp_mux_70_ comp_mux_00_ comp_mux_26_ vdd_d vss_d comp_mux_27_ / CKND2D1LVT
XXcomp_mux_72_ net2690 net2580 vdd_d vss_d comp_mux_29_ / CKND2D1LVT
XXcomp_mux_78_ comp_mux_34_ comp_mux_04_ vdd_d vss_d comp_mux_35_ / CKND2D1LVT
XXcomp_mux_76_ net2581 net2738 vdd_d vss_d comp_mux_33_ / CKND2D2LVT
XXcomp_mux_83_ comp_mux_35_ comp_mux_39_ spi_bits[178] vdd_d vss_d 
+ comp_mux_40_ / ND3D2LVT
XXcomp_mux_85_ comp_mux_31_ comp_mux_40_ net2467 vdd_d vss_d comp_mux_42_ / 
+ ND3D2LVT
XXspi_reg_0_ net2 vdd_d vss_d spi_reg_enable / CKND1LVT
XXclkbuf_0_seq_init net2807 vdd_d vss_d clknet_0_seq_init / BUFFD16LVT
XXclkbuf_4_15_f_spi_sclk clknet_3_7_0_spi_sclk vdd_d vss_d 
+ clknet_4_15_leaf_spi_sclk / BUFFD16LVT
XXclkload5 clknet_4_11_leaf_spi_sclk vdd_d vss_d _unconnected_186 / BUFFD16LVT
XXclkbuf_4_0_f_spi_sclk clknet_3_0_0_spi_sclk vdd_d vss_d 
+ clknet_4_0_leaf_spi_sclk / BUFFD16LVT
XXclkbuf_3_5_0_spi_sclk clknet_0_spi_sclk vdd_d vss_d clknet_3_5_0_spi_sclk / 
+ BUFFD16LVT
XXclkbuf_4_1_f_spi_sclk clknet_3_0_0_spi_sclk vdd_d vss_d 
+ clknet_4_1_leaf_spi_sclk / BUFFD16LVT
XXclkbuf_3_6_0_spi_sclk net2870 vdd_d vss_d clknet_3_6_0_spi_sclk / BUFFD16LVT
XXclkbuf_4_4_f_spi_sclk clknet_3_2_0_spi_sclk vdd_d vss_d 
+ clknet_4_4_leaf_spi_sclk / BUFFD16LVT
XXclkbuf_3_7_0_spi_sclk net2870 vdd_d vss_d clknet_3_7_0_spi_sclk / BUFFD16LVT
XXclkbuf_4_3_f_spi_sclk clknet_3_1_0_spi_sclk vdd_d vss_d 
+ clknet_4_3_leaf_spi_sclk / BUFFD16LVT
XXclkbuf_4_2_f_spi_sclk clknet_3_1_0_spi_sclk vdd_d vss_d 
+ clknet_4_2_leaf_spi_sclk / BUFFD16LVT
XXclkbuf_4_8_f_spi_sclk clknet_3_4_0_spi_sclk vdd_d vss_d 
+ clknet_4_8_leaf_spi_sclk / BUFFD16LVT
XXclkbuf_4_7_f_spi_sclk clknet_3_3_0_spi_sclk vdd_d vss_d 
+ clknet_4_7_leaf_spi_sclk / BUFFD16LVT
XXclkbuf_4_14_f_spi_sclk clknet_3_7_0_spi_sclk vdd_d vss_d 
+ clknet_4_14_leaf_spi_sclk / BUFFD16LVT
XXclkbuf_4_12_f_spi_sclk clknet_3_6_0_spi_sclk vdd_d vss_d 
+ clknet_4_12_leaf_spi_sclk / BUFFD16LVT
XXclkbuf_4_6_f_spi_sclk clknet_3_3_0_spi_sclk vdd_d vss_d 
+ clknet_4_6_leaf_spi_sclk / BUFFD16LVT
XXclkbuf_4_5_f_spi_sclk clknet_3_2_0_spi_sclk vdd_d vss_d 
+ clknet_4_5_leaf_spi_sclk / BUFFD16LVT
XXclkbuf_4_11_f_spi_sclk clknet_3_5_0_spi_sclk vdd_d vss_d 
+ clknet_4_11_leaf_spi_sclk / BUFFD16LVT
XXclkbuf_4_10_f_spi_sclk clknet_3_5_0_spi_sclk vdd_d vss_d 
+ clknet_4_10_leaf_spi_sclk / BUFFD16LVT
XXclkbuf_4_9_f_spi_sclk clknet_3_4_0_spi_sclk vdd_d vss_d 
+ clknet_4_9_leaf_spi_sclk / BUFFD16LVT
XXclkbuf_3_1_0_spi_sclk net2871 vdd_d vss_d clknet_3_1_0_spi_sclk / BUFFD16LVT
XXclkbuf_3_4_0_spi_sclk clknet_0_spi_sclk vdd_d vss_d clknet_3_4_0_spi_sclk / 
+ BUFFD16LVT
XXclkbuf_3_3_0_spi_sclk net2869 vdd_d vss_d clknet_3_3_0_spi_sclk / BUFFD16LVT
XXclkbuf_3_2_0_spi_sclk net2869 vdd_d vss_d clknet_3_2_0_spi_sclk / BUFFD16LVT
XXclkbuf_3_0_0_spi_sclk net2871 vdd_d vss_d clknet_3_0_0_spi_sclk / BUFFD16LVT
XXclkbuf_1_0_f_seq_logic clknet_0_seq_logic vdd_d vss_d 
+ clknet_1_0_leaf_seq_logic / BUFFD16LVT
XXclkbuf_0_seq_logic net2851 vdd_d vss_d clknet_0_seq_logic / BUFFD16LVT
XXclkbuf_0_spi_sclk net2867 vdd_d vss_d clknet_0_spi_sclk / BUFFD16LVT
XXclkbuf_1_1_f_seq_logic clknet_0_seq_logic vdd_d vss_d 
+ clknet_1_1_leaf_seq_logic / BUFFD16LVT
XXclkbuf_1_0_f_seq_comp clknet_0_seq_comp vdd_d vss_d clknet_1_0_leaf_seq_comp 
+ / BUFFD16LVT
XXclkbuf_1_1_f_seq_comp clknet_0_seq_comp vdd_d vss_d clknet_1_1_leaf_seq_comp 
+ / BUFFD16LVT
XXclkbuf_1_0_f_seq_samp clknet_0_seq_samp vdd_d vss_d clknet_1_0_leaf_seq_samp 
+ / BUFFD16LVT
XXclkbuf_0_seq_samp net2821 vdd_d vss_d clknet_0_seq_samp / BUFFD16LVT
XXclkbuf_1_0_f_seq_init clknet_0_seq_init vdd_d vss_d clknet_1_0_leaf_seq_init 
+ / BUFFD16LVT
XXclkbuf_1_1_f_seq_init clknet_0_seq_init vdd_d vss_d clknet_1_1_leaf_seq_init 
+ / BUFFD16LVT
XXclkbuf_1_1_f_seq_samp clknet_0_seq_samp vdd_d vss_d clknet_1_1_leaf_seq_samp 
+ / BUFFD16LVT
XXclkbuf_0_seq_comp net2837 vdd_d vss_d clknet_0_seq_comp / BUFFD16LVT
XXclkbuf_4_13_f_spi_sclk clknet_3_6_0_spi_sclk vdd_d vss_d 
+ clknet_4_13_leaf_spi_sclk / BUFFD16LVT
XXspi_reg_sdo_dff_dffe net2725 net2806 spi_bits[179] net2689 net5 
+ _unconnected_0 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[0] net2706 clknet_4_7_leaf_spi_sclk net3 
+ net2889 spi_bits[0] _unconnected_1 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[100] net2708 clknet_4_6_leaf_spi_sclk 
+ spi_bits[99] net2675 spi_bits[100] _unconnected_2 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[101] net2708 clknet_4_0_leaf_spi_sclk 
+ spi_bits[100] net2675 spi_bits[101] _unconnected_3 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[102] net2708 clknet_4_0_leaf_spi_sclk 
+ spi_bits[101] net2675 spi_bits[102] _unconnected_4 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[103] net2708 clknet_4_0_leaf_spi_sclk 
+ spi_bits[102] net2675 spi_bits[103] _unconnected_5 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[104] net2708 clknet_4_0_leaf_spi_sclk 
+ spi_bits[103] net2675 spi_bits[104] _unconnected_6 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[105] net2725 clknet_4_0_leaf_spi_sclk 
+ spi_bits[104] net2689 spi_bits[105] _unconnected_7 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[106] net2712 clknet_4_8_leaf_spi_sclk 
+ spi_bits[105] net2678 spi_bits[106] _unconnected_8 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[107] net2717 clknet_4_10_leaf_spi_sclk 
+ spi_bits[106] net2682 spi_bits[107] _unconnected_9 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[108] net2717 clknet_4_10_leaf_spi_sclk 
+ spi_bits[107] net2682 spi_bits[108] _unconnected_10 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[109] net2717 clknet_4_10_leaf_spi_sclk 
+ spi_bits[108] net2682 spi_bits[109] _unconnected_11 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[10] net2720 clknet_4_10_leaf_spi_sclk 
+ spi_bits[9] net2684 spi_bits[10] _unconnected_12 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[110] net2719 clknet_4_11_leaf_spi_sclk 
+ spi_bits[109] net2684 spi_bits[110] _unconnected_13 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[111] net2719 clknet_4_11_leaf_spi_sclk 
+ spi_bits[110] net2684 spi_bits[111] _unconnected_14 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[112] net2720 clknet_4_10_leaf_spi_sclk 
+ spi_bits[111] net2684 spi_bits[112] _unconnected_15 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[113] net2721 clknet_4_12_leaf_spi_sclk 
+ spi_bits[112] net2685 spi_bits[113] _unconnected_16 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[114] net2723 clknet_4_12_leaf_spi_sclk 
+ spi_bits[113] net2687 spi_bits[114] _unconnected_17 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[115] net2723 clknet_4_14_leaf_spi_sclk 
+ spi_bits[114] net2687 spi_bits[115] _unconnected_18 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[116] net2723 clknet_4_14_leaf_spi_sclk 
+ spi_bits[115] net2687 spi_bits[116] _unconnected_19 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[117] net2723 clknet_4_14_leaf_spi_sclk 
+ spi_bits[116] net2687 spi_bits[117] _unconnected_20 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[118] net2723 clknet_4_14_leaf_spi_sclk 
+ spi_bits[117] net2687 spi_bits[118] _unconnected_21 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[119] net2723 clknet_4_14_leaf_spi_sclk 
+ spi_bits[118] net2687 spi_bits[119] _unconnected_22 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[11] net2716 clknet_4_10_leaf_spi_sclk 
+ spi_bits[10] net2682 spi_bits[11] _unconnected_23 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[120] net2711 clknet_4_2_leaf_spi_sclk 
+ net2635 net2677 spi_bits[120] _unconnected_24 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[121] net2694 clknet_4_4_leaf_spi_sclk 
+ net2630 net2662 spi_bits[121] _unconnected_25 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[122] net1 clknet_4_4_leaf_spi_sclk 
+ spi_bits[121] net2663 spi_bits[122] _unconnected_26 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[123] net1 clknet_4_4_leaf_spi_sclk 
+ spi_bits[122] net2663 spi_bits[123] _unconnected_27 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[124] net2692 clknet_4_4_leaf_spi_sclk 
+ spi_bits[123] net2663 spi_bits[124] _unconnected_28 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[125] net2692 clknet_4_4_leaf_spi_sclk 
+ spi_bits[124] net2663 spi_bits[125] _unconnected_29 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[126] net2692 clknet_4_4_leaf_spi_sclk 
+ spi_bits[125] net2663 spi_bits[126] _unconnected_30 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[127] net2695 clknet_4_4_leaf_spi_sclk 
+ spi_bits[126] net2664 spi_bits[127] _unconnected_31 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[128] net2724 clknet_4_1_leaf_spi_sclk 
+ net2622 net2688 spi_bits[128] _unconnected_32 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[129] net2724 clknet_4_1_leaf_spi_sclk 
+ spi_bits[128] net2688 spi_bits[129] _unconnected_33 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[12] net2717 clknet_4_10_leaf_spi_sclk 
+ spi_bits[11] net2682 spi_bits[12] _unconnected_34 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[130] net2724 clknet_4_1_leaf_spi_sclk 
+ spi_bits[129] net2688 spi_bits[130] _unconnected_35 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[131] net2709 clknet_4_1_leaf_spi_sclk 
+ spi_bits[130] net2688 spi_bits[131] _unconnected_36 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[132] net2709 clknet_4_1_leaf_spi_sclk 
+ spi_bits[131] net2676 spi_bits[132] _unconnected_37 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[133] net2725 clknet_4_0_leaf_spi_sclk 
+ spi_bits[132] net2689 spi_bits[133] _unconnected_38 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[134] net2712 clknet_4_2_leaf_spi_sclk 
+ spi_bits[133] net2678 spi_bits[134] _unconnected_39 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[135] net2713 clknet_4_9_leaf_spi_sclk 
+ spi_bits[134] net2679 spi_bits[135] _unconnected_40 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[136] net2713 clknet_4_8_leaf_spi_sclk 
+ spi_bits[135] net2679 spi_bits[136] _unconnected_41 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[137] net2713 clknet_4_8_leaf_spi_sclk 
+ spi_bits[136] net2679 spi_bits[137] _unconnected_42 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[138] net2713 clknet_4_8_leaf_spi_sclk 
+ spi_bits[137] net2680 spi_bits[138] _unconnected_43 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[139] net2714 clknet_4_8_leaf_spi_sclk 
+ spi_bits[138] net2680 spi_bits[139] _unconnected_44 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[13] net2717 clknet_4_10_leaf_spi_sclk 
+ spi_bits[12] net2682 spi_bits[13] _unconnected_45 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[140] net2714 clknet_4_8_leaf_spi_sclk 
+ spi_bits[139] net2680 spi_bits[140] _unconnected_46 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[141] net2714 clknet_4_8_leaf_spi_sclk 
+ spi_bits[140] net2680 spi_bits[141] _unconnected_47 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[142] net2722 clknet_4_12_leaf_spi_sclk 
+ spi_bits[141] net2686 spi_bits[142] _unconnected_48 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[143] net2722 clknet_4_14_leaf_spi_sclk 
+ spi_bits[142] net2686 spi_bits[143] _unconnected_49 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[144] net2722 clknet_4_14_leaf_spi_sclk 
+ spi_bits[143] net2686 spi_bits[144] _unconnected_50 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[145] net2722 clknet_4_14_leaf_spi_sclk 
+ spi_bits[144] net2686 spi_bits[145] _unconnected_51 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[146] net2722 clknet_4_14_leaf_spi_sclk 
+ spi_bits[145] net2686 spi_bits[146] _unconnected_52 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[147] net2722 clknet_4_12_leaf_spi_sclk 
+ spi_bits[146] net2686 spi_bits[147] _unconnected_53 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[148] net2725 clknet_4_1_leaf_spi_sclk 
+ net2599 net2689 spi_bits[148] _unconnected_54 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[149] net2698 clknet_4_4_leaf_spi_sclk 
+ net2596 net2667 spi_bits[149] _unconnected_55 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[14] net2717 clknet_4_10_leaf_spi_sclk 
+ spi_bits[13] net2682 spi_bits[14] _unconnected_56 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[150] net2699 clknet_4_4_leaf_spi_sclk 
+ spi_bits[149] net2771 spi_bits[150] _unconnected_57 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[151] net2768 clknet_4_4_leaf_spi_sclk 
+ net2782 net2771 spi_bits[151] _unconnected_58 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[152] net2875 clknet_4_5_leaf_spi_sclk 
+ net2781 net2874 spi_bits[152] _unconnected_59 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[153] net2875 clknet_4_5_leaf_spi_sclk 
+ spi_bits[152] net2874 spi_bits[153] _unconnected_60 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[154] net2875 clknet_4_5_leaf_spi_sclk 
+ spi_bits[153] net2874 spi_bits[154] _unconnected_61 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[155] net2700 clknet_4_4_leaf_spi_sclk 
+ net2779 net2667 spi_bits[155] _unconnected_62 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[156] net2700 clknet_4_6_leaf_spi_sclk 
+ net2778 net2669 spi_bits[156] _unconnected_63 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[157] net2766 clknet_4_0_leaf_spi_sclk 
+ net2774 net2669 spi_bits[157] _unconnected_64 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[158] net2766 clknet_4_0_leaf_spi_sclk 
+ net2884 net2769 spi_bits[158] _unconnected_65 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[159] net2765 clknet_4_7_leaf_spi_sclk 
+ net2773 net2670 spi_bits[159] _unconnected_66 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[160] net2765 clknet_4_7_leaf_spi_sclk 
+ net2876 net2670 spi_bits[160] _unconnected_68 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[161] net2765 clknet_4_1_leaf_spi_sclk 
+ spi_bits[160] net2670 spi_bits[161] _unconnected_69 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[162] net2702 clknet_4_3_leaf_spi_sclk 
+ net2882 net2670 spi_bits[162] _unconnected_70 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[163] net2702 clknet_4_9_leaf_spi_sclk 
+ spi_bits[162] net2671 spi_bits[163] _unconnected_71 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[164] net2703 clknet_4_9_leaf_spi_sclk 
+ spi_bits[163] net2671 spi_bits[164] _unconnected_72 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[165] net2703 clknet_4_11_leaf_spi_sclk 
+ net2885 net2671 spi_bits[165] _unconnected_73 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[166] net2703 clknet_4_11_leaf_spi_sclk 
+ spi_bits[165] net2672 spi_bits[166] _unconnected_74 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[167] net2703 clknet_4_11_leaf_spi_sclk 
+ spi_bits[166] net2672 spi_bits[167] _unconnected_75 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[168] net2704 clknet_4_13_leaf_spi_sclk 
+ spi_bits[167] net2672 spi_bits[168] _unconnected_76 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[169] net2704 clknet_4_13_leaf_spi_sclk 
+ spi_bits[168] net2672 spi_bits[169] _unconnected_77 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[16] net2719 clknet_4_11_leaf_spi_sclk 
+ spi_bits[15] net2683 spi_bits[16] _unconnected_78 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[170] net2704 clknet_4_15_leaf_spi_sclk 
+ spi_bits[169] net2673 spi_bits[170] _unconnected_79 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[171] net2705 clknet_4_15_leaf_spi_sclk 
+ spi_bits[170] net2673 spi_bits[171] _unconnected_80 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[172] net2705 clknet_4_15_leaf_spi_sclk 
+ spi_bits[171] net2673 spi_bits[172] _unconnected_81 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[173] net2763 clknet_4_15_leaf_spi_sclk 
+ spi_bits[172] net2764 spi_bits[173] _unconnected_82 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[174] net2763 clknet_4_14_leaf_spi_sclk 
+ spi_bits[173] net2764 spi_bits[174] _unconnected_83 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[175] net2763 clknet_4_15_leaf_spi_sclk 
+ spi_bits[174] net2764 spi_bits[175] _unconnected_84 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[176] net2721 clknet_4_12_leaf_spi_sclk 
+ net2586 net2685 spi_bits[176] _unconnected_85 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[177] net2712 clknet_4_2_leaf_spi_sclk 
+ net2582 net2678 spi_bits[177] _unconnected_86 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[178] net2712 clknet_4_2_leaf_spi_sclk 
+ spi_bits[177] net2678 spi_bits[178] _unconnected_87 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[179] net2711 clknet_4_2_leaf_spi_sclk 
+ spi_bits[178] net2678 spi_bits[179] _unconnected_88 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[17] net2718 clknet_4_8_leaf_spi_sclk 
+ spi_bits[16] net2683 spi_bits[17] _unconnected_89 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[18] net2718 clknet_4_9_leaf_spi_sclk 
+ spi_bits[17] net2681 spi_bits[18] _unconnected_90 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[19] net2718 clknet_4_8_leaf_spi_sclk 
+ spi_bits[18] net2681 spi_bits[19] _unconnected_91 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[1] net2716 clknet_4_2_leaf_spi_sclk 
+ net2659 net2681 spi_bits[1] _unconnected_92 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[20] net2716 clknet_4_9_leaf_spi_sclk 
+ spi_bits[19] net2681 spi_bits[20] _unconnected_93 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[21] net2717 clknet_4_11_leaf_spi_sclk 
+ spi_bits[20] net2682 spi_bits[21] _unconnected_94 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[22] net2718 clknet_4_8_leaf_spi_sclk 
+ spi_bits[21] net2683 spi_bits[22] _unconnected_95 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[23] net2718 clknet_4_10_leaf_spi_sclk 
+ spi_bits[22] net2683 spi_bits[23] _unconnected_96 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[24] net2716 clknet_4_9_leaf_spi_sclk 
+ spi_bits[23] net2681 spi_bits[24] _unconnected_97 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[25] net2718 clknet_4_8_leaf_spi_sclk 
+ spi_bits[24] net2681 spi_bits[25] _unconnected_98 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[26] net2718 clknet_4_8_leaf_spi_sclk 
+ spi_bits[25] net2683 spi_bits[26] _unconnected_99 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[27] net2720 clknet_4_12_leaf_spi_sclk 
+ net2873 net2684 spi_bits[27] _unconnected_100 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[28] net2720 clknet_4_13_leaf_spi_sclk 
+ spi_bits[27] net2684 spi_bits[28] _unconnected_101 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[29] net2719 clknet_4_13_leaf_spi_sclk 
+ spi_bits[28] net2684 spi_bits[29] _unconnected_102 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[2] net2718 clknet_4_8_leaf_spi_sclk 
+ spi_bits[1] net2683 spi_bits[2] _unconnected_103 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[30] net2716 clknet_4_11_leaf_spi_sclk 
+ spi_bits[29] net2682 spi_bits[30] _unconnected_104 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[31] net2712 clknet_4_2_leaf_spi_sclk 
+ spi_bits[30] net2678 spi_bits[31] _unconnected_105 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[32] net2712 clknet_4_2_leaf_spi_sclk 
+ spi_bits[31] net2678 spi_bits[32] _unconnected_106 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[33] net2711 clknet_4_2_leaf_spi_sclk 
+ spi_bits[32] net2677 spi_bits[33] _unconnected_107 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[34] net2711 clknet_4_2_leaf_spi_sclk 
+ spi_bits[33] net2677 spi_bits[34] _unconnected_108 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[35] net2708 clknet_4_6_leaf_spi_sclk 
+ spi_bits[34] net2675 spi_bits[35] _unconnected_109 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[36] net2708 clknet_4_6_leaf_spi_sclk 
+ spi_bits[35] net2675 spi_bits[36] _unconnected_110 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[37] net2708 clknet_4_6_leaf_spi_sclk 
+ spi_bits[36] net2675 spi_bits[37] _unconnected_111 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[38] net2708 clknet_4_6_leaf_spi_sclk 
+ spi_bits[37] net2675 spi_bits[38] _unconnected_112 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[39] net2711 clknet_4_1_leaf_spi_sclk 
+ spi_bits[38] net2677 spi_bits[39] _unconnected_113 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[3] net2720 clknet_4_10_leaf_spi_sclk 
+ spi_bits[2] net2684 spi_bits[3] _unconnected_114 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[40] net2711 clknet_4_2_leaf_spi_sclk 
+ spi_bits[39] net2677 spi_bits[40] _unconnected_115 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[41] net2708 clknet_4_0_leaf_spi_sclk 
+ spi_bits[40] net2675 spi_bits[41] _unconnected_116 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[42] net2707 clknet_4_0_leaf_spi_sclk 
+ spi_bits[41] net2689 spi_bits[42] _unconnected_117 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[43] net2710 clknet_4_1_leaf_spi_sclk 
+ spi_bits[42] net2677 spi_bits[43] _unconnected_118 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[44] net2710 clknet_4_1_leaf_spi_sclk 
+ spi_bits[43] net2677 spi_bits[44] _unconnected_119 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[45] net2715 clknet_4_3_leaf_spi_sclk 
+ spi_bits[44] net2676 spi_bits[45] _unconnected_120 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[46] net2710 clknet_4_1_leaf_spi_sclk 
+ spi_bits[45] net2677 spi_bits[46] _unconnected_121 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[47] net2707 clknet_4_1_leaf_spi_sclk 
+ spi_bits[46] net2674 spi_bits[47] _unconnected_122 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[48] net2725 clknet_4_1_leaf_spi_sclk 
+ spi_bits[47] net2689 spi_bits[48] _unconnected_123 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[49] net2711 clknet_4_3_leaf_spi_sclk 
+ spi_bits[48] net2677 spi_bits[49] _unconnected_124 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[4] net2720 clknet_4_12_leaf_spi_sclk 
+ net2872 net2684 spi_bits[4] _unconnected_125 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[50] net2711 clknet_4_2_leaf_spi_sclk 
+ spi_bits[49] net2677 spi_bits[50] _unconnected_126 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[51] net2725 clknet_4_1_leaf_spi_sclk 
+ spi_bits[50] net2689 spi_bits[51] _unconnected_127 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[52] net2707 clknet_4_1_leaf_spi_sclk 
+ spi_bits[51] net2689 spi_bits[52] _unconnected_128 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[53] net2715 clknet_4_3_leaf_spi_sclk 
+ spi_bits[52] net2676 spi_bits[53] _unconnected_129 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[54] net2715 clknet_4_3_leaf_spi_sclk 
+ spi_bits[53] net2676 spi_bits[54] _unconnected_130 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[55] net2707 clknet_4_0_leaf_spi_sclk 
+ spi_bits[54] net2674 spi_bits[55] _unconnected_131 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[56] net2710 clknet_4_1_leaf_spi_sclk 
+ spi_bits[55] net2677 spi_bits[56] _unconnected_132 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[57] net2715 clknet_4_3_leaf_spi_sclk 
+ spi_bits[56] net2681 spi_bits[57] _unconnected_133 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[58] net2715 clknet_4_1_leaf_spi_sclk 
+ spi_bits[57] net2676 spi_bits[58] _unconnected_134 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[59] net2715 clknet_4_3_leaf_spi_sclk 
+ spi_bits[58] net2681 spi_bits[59] _unconnected_135 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[5] net2720 clknet_4_13_leaf_spi_sclk 
+ spi_bits[4] net2684 spi_bits[5] _unconnected_136 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[60] net2715 clknet_4_3_leaf_spi_sclk 
+ spi_bits[59] net2676 spi_bits[60] _unconnected_137 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[61] net2710 clknet_4_3_leaf_spi_sclk 
+ spi_bits[60] net2676 spi_bits[61] _unconnected_138 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[62] net2706 clknet_4_7_leaf_spi_sclk 
+ spi_bits[61] net2889 spi_bits[62] _unconnected_139 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[63] net2706 clknet_4_7_leaf_spi_sclk 
+ spi_bits[62] net2889 spi_bits[63] _unconnected_140 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[64] net2693 clknet_4_5_leaf_spi_sclk 
+ spi_bits[63] net2661 spi_bits[64] _unconnected_141 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[65] net2692 clknet_4_5_leaf_spi_sclk 
+ spi_bits[64] net2663 spi_bits[65] _unconnected_142 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[66] net2692 clknet_4_5_leaf_spi_sclk 
+ spi_bits[65] net2663 spi_bits[66] _unconnected_143 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[67] net2692 clknet_4_5_leaf_spi_sclk 
+ spi_bits[66] net2663 spi_bits[67] _unconnected_144 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[68] net2692 clknet_4_5_leaf_spi_sclk 
+ spi_bits[67] net2663 spi_bits[68] _unconnected_145 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[69] net2692 clknet_4_4_leaf_spi_sclk 
+ spi_bits[68] net2663 spi_bits[69] _unconnected_146 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[6] net2717 clknet_4_10_leaf_spi_sclk 
+ spi_bits[5] net2682 spi_bits[6] _unconnected_147 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[70] net2692 clknet_4_5_leaf_spi_sclk 
+ spi_bits[69] net2663 spi_bits[70] _unconnected_148 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[71] net2693 clknet_4_7_leaf_spi_sclk 
+ spi_bits[70] net2889 spi_bits[71] _unconnected_149 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[72] net2706 clknet_4_6_leaf_spi_sclk 
+ spi_bits[71] net2674 spi_bits[72] _unconnected_150 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[73] net2707 clknet_4_0_leaf_spi_sclk 
+ spi_bits[72] net2674 spi_bits[73] _unconnected_151 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[74] net2707 clknet_4_0_leaf_spi_sclk 
+ spi_bits[73] net2674 spi_bits[74] _unconnected_152 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[75] net2709 clknet_4_1_leaf_spi_sclk 
+ spi_bits[74] net2676 spi_bits[75] _unconnected_153 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[76] net2709 clknet_4_1_leaf_spi_sclk 
+ spi_bits[75] net2676 spi_bits[76] _unconnected_154 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[77] net2710 clknet_4_1_leaf_spi_sclk 
+ spi_bits[76] net2676 spi_bits[77] _unconnected_155 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[78] net2716 clknet_4_9_leaf_spi_sclk 
+ spi_bits[77] net2681 spi_bits[78] _unconnected_156 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[79] net2718 clknet_4_10_leaf_spi_sclk 
+ spi_bits[78] net2683 spi_bits[79] _unconnected_157 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[7] net2717 clknet_4_11_leaf_spi_sclk 
+ spi_bits[6] net2682 spi_bits[7] _unconnected_158 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[80] net2719 clknet_4_10_leaf_spi_sclk 
+ spi_bits[79] net2683 spi_bits[80] _unconnected_159 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[81] net2719 clknet_4_11_leaf_spi_sclk 
+ spi_bits[80] net2683 spi_bits[81] _unconnected_160 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[82] net2719 clknet_4_11_leaf_spi_sclk 
+ spi_bits[81] net2683 spi_bits[82] _unconnected_161 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[83] net2719 clknet_4_10_leaf_spi_sclk 
+ spi_bits[82] net2683 spi_bits[83] _unconnected_162 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[84] net2719 clknet_4_11_leaf_spi_sclk 
+ spi_bits[83] net2683 spi_bits[84] _unconnected_163 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[85] net2720 clknet_4_13_leaf_spi_sclk 
+ spi_bits[84] net2685 spi_bits[85] _unconnected_164 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[86] net2723 clknet_4_12_leaf_spi_sclk 
+ spi_bits[85] net2687 spi_bits[86] _unconnected_165 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[87] net2723 clknet_4_14_leaf_spi_sclk 
+ spi_bits[86] net2687 spi_bits[87] _unconnected_166 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[88] net2723 clknet_4_15_leaf_spi_sclk 
+ spi_bits[87] net2687 spi_bits[88] _unconnected_167 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[89] net2723 clknet_4_15_leaf_spi_sclk 
+ spi_bits[88] net2687 spi_bits[89] _unconnected_168 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[8] net2719 clknet_4_10_leaf_spi_sclk 
+ spi_bits[7] net2684 spi_bits[8] _unconnected_169 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[90] net2723 clknet_4_15_leaf_spi_sclk 
+ spi_bits[89] net2687 spi_bits[90] _unconnected_170 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[91] net2723 clknet_4_14_leaf_spi_sclk 
+ spi_bits[90] net2687 spi_bits[91] _unconnected_171 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[92] net2716 clknet_4_9_leaf_spi_sclk 
+ net2480 net2681 spi_bits[92] _unconnected_172 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[93] net2693 clknet_4_7_leaf_spi_sclk 
+ net2477 net2661 spi_bits[93] _unconnected_173 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[94] net2693 clknet_4_5_leaf_spi_sclk 
+ spi_bits[93] net2661 spi_bits[94] _unconnected_174 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[95] net2693 clknet_4_5_leaf_spi_sclk 
+ spi_bits[94] net2663 spi_bits[95] _unconnected_175 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[96] net2693 clknet_4_4_leaf_spi_sclk 
+ spi_bits[95] net2663 spi_bits[96] _unconnected_176 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[97] net2692 clknet_4_4_leaf_spi_sclk 
+ spi_bits[96] net2663 spi_bits[97] _unconnected_177 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[98] net2693 clknet_4_7_leaf_spi_sclk 
+ spi_bits[97] net2663 spi_bits[98] _unconnected_178 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[99] net2693 clknet_4_7_leaf_spi_sclk 
+ spi_bits[98] net2889 spi_bits[99] _unconnected_179 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[9] net2719 clknet_4_10_leaf_spi_sclk 
+ spi_bits[8] net2684 spi_bits[9] _unconnected_180 vdd_d vss_d / EDFCND2LVT
XXspi_reg_shift_stage_dff_inst_dffe[15] net2720 clknet_4_10_leaf_spi_sclk 
+ spi_bits[14] net2684 spi_bits[15] _unconnected_67 vdd_d vss_d / EDFCND4LVT
XXplace2467 comp_mux_41_ vdd_d vss_d net2467 / CKBD2LVT
XXplace2480 net2479 vdd_d vss_d net2480 / CKBD2LVT
XXplace2478 net2477 vdd_d vss_d net2478 / CKBD2LVT
XXplace2516 spi_bits[4] vdd_d vss_d net2516 / CKBD2LVT
XXplace2518 net2516 vdd_d vss_d net2518 / CKBD2LVT
XXplace2590 net2775 vdd_d vss_d net2590 / CKBD2LVT
XXplace2597 net2596 vdd_d vss_d net2597 / CKBD2LVT
XXplace2600 spi_bits[147] vdd_d vss_d net2600 / CKBD2LVT
XXplace2599 net2598 vdd_d vss_d net2599 / CKBD2LVT
XXplace2607 spi_bits[140] vdd_d vss_d net2607 / CKBD2LVT
XXplace2615 spi_bits[133] vdd_d vss_d net2615 / CKBD2LVT
XXplace2609 spi_bits[139] vdd_d vss_d net2609 / CKBD2LVT
XXplace2631 net2630 vdd_d vss_d net2631 / CKBD2LVT
XXplace2620 spi_bits[129] vdd_d vss_d net2620 / CKBD2LVT
XXplace2582 net2881 vdd_d vss_d net2582 / CKBD2LVT
XXplace2580 net2881 vdd_d vss_d net2580 / CKBD2LVT
XXplace2581 net2580 vdd_d vss_d net2581 / CKBD2LVT
XXplace2579 spi_bits[176] vdd_d vss_d net2579 / CKBD2LVT
XXplace2586 net2585 vdd_d vss_d net2586 / CKBD2LVT
XXplace2636 spi_bits[119] vdd_d vss_d net2636 / CKBD2LVT
XXplace2644 spi_bits[111] vdd_d vss_d net2644 / CKBD2LVT
XXplace2643 spi_bits[112] vdd_d vss_d net2643 / CKBD2LVT
XXplace2635 net2634 vdd_d vss_d net2635 / CKBD2LVT
XXplace2642 spi_bits[113] vdd_d vss_d net2642 / CKBD2LVT
XXplace2686 net2685 vdd_d vss_d net2686 / CKBD2LVT
XXplace2687 net2685 vdd_d vss_d net2687 / CKBD2LVT
XXplace2688 net2676 vdd_d vss_d net2688 / CKBD2LVT
XXplace2689 net2674 vdd_d vss_d net2689 / CKBD2LVT
XXplace2645 spi_bits[110] vdd_d vss_d net2645 / CKBD2LVT
XXplace2654 spi_bits[102] vdd_d vss_d net2654 / CKBD2LVT
XXplace2653 spi_bits[103] vdd_d vss_d net2653 / CKBD2LVT
XXplace2648 spi_bits[108] vdd_d vss_d net2648 / CKBD2LVT
XXplace2652 spi_bits[104] vdd_d vss_d net2652 / CKBD2LVT
XXplace2651 spi_bits[105] vdd_d vss_d net2651 / CKBD2LVT
XXplace2649 spi_bits[107] vdd_d vss_d net2649 / CKBD2LVT
XXplace2650 spi_bits[106] vdd_d vss_d net2650 / CKBD2LVT
XXplace2655 spi_bits[101] vdd_d vss_d net2655 / CKBD2LVT
XXplace2656 spi_bits[100] vdd_d vss_d net2656 / CKBD2LVT
XXplace2685 net2684 vdd_d vss_d net2685 / CKBD2LVT
XXplace2647 spi_bits[109] vdd_d vss_d net2647 / CKBD2LVT
XXplace2601 spi_bits[146] vdd_d vss_d net2601 / CKBD2LVT
XXplace2663 net2662 vdd_d vss_d net2663 / CKBD2LVT
XXplace2661 spi_reg_enable vdd_d vss_d net2661 / CKBD2LVT
XXplace2662 net2661 vdd_d vss_d net2662 / CKBD2LVT
XXplace2701 net2700 vdd_d vss_d net2701 / CKBD2LVT
XXplace2699 net2698 vdd_d vss_d net2699 / CKBD2LVT
XXplace2700 net2698 vdd_d vss_d net2700 / CKBD2LVT
XXplace2690 comp_mux_28_ vdd_d vss_d net2690 / CKBD2LVT
XXplace2703 net2702 vdd_d vss_d net2703 / CKBD2LVT
XXplace2698 net2697 vdd_d vss_d net2698 / CKBD2LVT
XXplace2705 net2704 vdd_d vss_d net2705 / CKBD2LVT
XXplace2721 net2720 vdd_d vss_d net2721 / CKBD2LVT
XXplace2695 net2694 vdd_d vss_d net2695 / CKBD2LVT
XXplace2711 net2710 vdd_d vss_d net2711 / CKBD2LVT
XXplace2713 net2712 vdd_d vss_d net2713 / CKBD2LVT
XXplace2710 net2709 vdd_d vss_d net2710 / CKBD2LVT
XXplace2709 net2707 vdd_d vss_d net2709 / CKBD2LVT
XXplace2719 net2718 vdd_d vss_d net2719 / CKBD2LVT
XXplace2706 net2693 vdd_d vss_d net2706 / CKBD2LVT
XXplace2707 net2706 vdd_d vss_d net2707 / CKBD2LVT
XXplace2702 net2765 vdd_d vss_d net2702 / CKBD2LVT
XXplace2704 net2703 vdd_d vss_d net2704 / CKBD2LVT
XXplace2658 spi_bits[0] vdd_d vss_d net2658 / CKBD2LVT
XXplace2677 net2676 vdd_d vss_d net2677 / CKBD2LVT
XXplace2684 net2683 vdd_d vss_d net2684 / CKBD2LVT
XXplace2659 net2658 vdd_d vss_d net2659 / CKBD2LVT
XXplace2712 net2711 vdd_d vss_d net2712 / CKBD2LVT
XXplace2714 net2713 vdd_d vss_d net2714 / CKBD2LVT
XXplace2676 net2674 vdd_d vss_d net2676 / CKBD2LVT
XXplace2722 net2721 vdd_d vss_d net2722 / CKBD2LVT
XXplace2675 net2674 vdd_d vss_d net2675 / CKBD2LVT
XXplace2720 net2719 vdd_d vss_d net2720 / CKBD2LVT
XXplace2717 net2716 vdd_d vss_d net2717 / CKBD2LVT
XXplace2718 net2716 vdd_d vss_d net2718 / CKBD2LVT
XXplace2716 net2715 vdd_d vss_d net2716 / CKBD2LVT
XXplace2715 net2710 vdd_d vss_d net2715 / CKBD2LVT
XXplace2683 net2681 vdd_d vss_d net2683 / CKBD2LVT
XXplace2682 net2681 vdd_d vss_d net2682 / CKBD2LVT
XXplace2681 net2676 vdd_d vss_d net2681 / CKBD2LVT
XXplace2680 net2679 vdd_d vss_d net2680 / CKBD2LVT
XXplace2660 net2659 vdd_d vss_d net2660 / CKBD2LVT
XXplace2679 net2678 vdd_d vss_d net2679 / CKBD2LVT
XXplace2678 net2677 vdd_d vss_d net2678 / CKBD2LVT
XXplace2723 net2721 vdd_d vss_d net2723 / CKBD2LVT
XXplace2725 net2707 vdd_d vss_d net2725 / CKBD2LVT
XXplace2724 net2709 vdd_d vss_d net2724 / CKBD2LVT
XXplace2694 net2693 vdd_d vss_d net2694 / CKBD2LVT
XXplace2693 net2692 vdd_d vss_d net2693 / CKBD2LVT
XXplace2692 net1 vdd_d vss_d net2692 / CKBD2LVT
XXplace2741 net2740 vdd_d vss_d net2741 / CKBD2LVT
XXplace2732 net2731 vdd_d vss_d net2732 / CKBD2LVT
XXplace2728 net2727 vdd_d vss_d net2728 / CKBD2LVT
XXplace2734 net2733 vdd_d vss_d net2734 / CKBD2LVT
XXwire1414 net2466 vdd_d vss_d spi_sdo / CKBD2LVT
XXplace2664 net2662 vdd_d vss_d net2664 / CKBD2LVT
XXplace2667 net2666 vdd_d vss_d net2667 / CKBD2LVT
XXplace2669 net2667 vdd_d vss_d net2669 / CKBD2LVT
XXplace2668 net2667 vdd_d vss_d net2668 / CKBD2LVT
XXplace2671 net2670 vdd_d vss_d net2671 / CKBD2LVT
XXplace2670 net2769 vdd_d vss_d net2670 / CKBD2LVT
XXplace2672 net2671 vdd_d vss_d net2672 / CKBD2LVT
XXplace2674 net2889 vdd_d vss_d net2674 / CKBD2LVT
XXplace2673 net2672 vdd_d vss_d net2673 / CKBD2LVT
XXplace2637 spi_bits[118] vdd_d vss_d net2637 / CKBD2LVT
XXplace2536 spi_bits[3] vdd_d vss_d net2536 / CKBD2LVT
XXplace2538 net2536 vdd_d vss_d net2538 / CKBD2LVT
XXplace2479 spi_bits[91] vdd_d vss_d net2479 / CKBD2LVT
XXplace2708 net2707 vdd_d vss_d net2708 / CKBD2LVT
XXplace2468 comp_mux_00_ vdd_d vss_d net2468 / CKBD2LVT
XXplace2487 spi_bits[63] vdd_d vss_d net2487 / CKBD2LVT
XXplace2489 spi_bits[63] vdd_d vss_d net2489 / CKBD2LVT
XXplace2484 spi_bits[71] vdd_d vss_d net2484 / CKBD2LVT
XXplace2476 spi_bits[93] vdd_d vss_d net2476 / CKBD2LVT
XXplace2472 spi_bits[97] vdd_d vss_d net2472 / CKBD2LVT
XXplace2471 spi_bits[98] vdd_d vss_d net2471 / CKBD2LVT
XXplace2470 spi_bits[99] vdd_d vss_d net2470 / CKBD2LVT
XXplace2473 spi_bits[96] vdd_d vss_d net2473 / CKBD2LVT
XXplace2474 spi_bits[95] vdd_d vss_d net2474 / CKBD2LVT
XXplace2475 spi_bits[94] vdd_d vss_d net2475 / CKBD2LVT
XXplace2602 spi_bits[145] vdd_d vss_d net2602 / CKBD2LVT
XXplace2603 spi_bits[144] vdd_d vss_d net2603 / CKBD2LVT
XXplace2604 spi_bits[143] vdd_d vss_d net2604 / CKBD2LVT
XXplace2605 spi_bits[142] vdd_d vss_d net2605 / CKBD2LVT
XXplace2606 spi_bits[141] vdd_d vss_d net2606 / CKBD2LVT
XXplace2610 spi_bits[138] vdd_d vss_d net2610 / CKBD2LVT
XXplace2611 spi_bits[137] vdd_d vss_d net2611 / CKBD2LVT
XXplace2612 spi_bits[136] vdd_d vss_d net2612 / CKBD2LVT
XXplace2613 spi_bits[135] vdd_d vss_d net2613 / CKBD2LVT
XXplace2614 spi_bits[134] vdd_d vss_d net2614 / CKBD2LVT
XXplace2616 spi_bits[132] vdd_d vss_d net2616 / CKBD2LVT
XXplace2617 spi_bits[131] vdd_d vss_d net2617 / CKBD2LVT
XXplace2618 spi_bits[130] vdd_d vss_d net2618 / CKBD2LVT
XXplace2621 spi_bits[128] vdd_d vss_d net2621 / CKBD2LVT
XXplace2623 net2622 vdd_d vss_d net2623 / CKBD2LVT
XXplace2624 spi_bits[126] vdd_d vss_d net2624 / CKBD2LVT
XXplace2625 spi_bits[125] vdd_d vss_d net2625 / CKBD2LVT
XXplace2626 spi_bits[124] vdd_d vss_d net2626 / CKBD2LVT
XXplace2627 spi_bits[123] vdd_d vss_d net2627 / CKBD2LVT
XXplace2628 spi_bits[122] vdd_d vss_d net2628 / CKBD2LVT
XXplace2629 spi_bits[121] vdd_d vss_d net2629 / CKBD2LVT
XXplace2638 spi_bits[117] vdd_d vss_d net2638 / CKBD2LVT
XXplace2639 spi_bits[116] vdd_d vss_d net2639 / CKBD2LVT
XXplace2640 spi_bits[115] vdd_d vss_d net2640 / CKBD2LVT
XXplace2641 spi_bits[114] vdd_d vss_d net2641 / CKBD2LVT
XXplace2745 net2744 vdd_d vss_d net2745 / CKBD2LVT
XXplace2738 net2737 vdd_d vss_d net2738 / CKBD2LVT
XXplace2736 net2735 vdd_d vss_d net2736 / CKBD2LVT
XXplace2749 net2748 vdd_d vss_d net2749 / CKBD2LVT
XXplace2752 net2751 vdd_d vss_d net2752 / CKBD2LVT
XXplace2756 net2755 vdd_d vss_d net2756 / CKBD2LVT
XXplace2759 net2758 vdd_d vss_d net2759 / CKBD2LVT
XXplace2762 net2761 vdd_d vss_d net2762 / CKBD2LVT
XXFILLER_20_320 vdd_d vss_d / DCAP64LVT
XXFILLER_20_256 vdd_d vss_d / DCAP64LVT
XXFILLER_20_64 vdd_d vss_d / DCAP64LVT
XXFILLER_20_0 vdd_d vss_d / DCAP64LVT
XXFILLER_17_808 vdd_d vss_d / DCAP64LVT
XXFILLER_16_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_16_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_16_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_16_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_16_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_16_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_16_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_16_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_19_1427 vdd_d vss_d / DCAP64LVT
XXFILLER_19_1555 vdd_d vss_d / DCAP64LVT
XXFILLER_19_1491 vdd_d vss_d / DCAP64LVT
XXFILLER_16_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_16_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_16_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_16_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_19_1299 vdd_d vss_d / DCAP64LVT
XXFILLER_16_832 vdd_d vss_d / DCAP64LVT
XXFILLER_16_896 vdd_d vss_d / DCAP64LVT
XXFILLER_16_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_16_960 vdd_d vss_d / DCAP64LVT
XXFILLER_16_768 vdd_d vss_d / DCAP64LVT
XXFILLER_16_704 vdd_d vss_d / DCAP64LVT
XXFILLER_16_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_16_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_16_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_16_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_16_576 vdd_d vss_d / DCAP64LVT
XXFILLER_16_640 vdd_d vss_d / DCAP64LVT
XXFILLER_16_0 vdd_d vss_d / DCAP64LVT
XXFILLER_16_128 vdd_d vss_d / DCAP64LVT
XXFILLER_16_64 vdd_d vss_d / DCAP64LVT
XXFILLER_16_256 vdd_d vss_d / DCAP64LVT
XXFILLER_16_192 vdd_d vss_d / DCAP64LVT
XXFILLER_16_384 vdd_d vss_d / DCAP64LVT
XXFILLER_16_320 vdd_d vss_d / DCAP64LVT
XXFILLER_15_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_15_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_15_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_15_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_15_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_15_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_15_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_18_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_15_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_15_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_15_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_15_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_15_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_15_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_15_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_15_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_15_512 vdd_d vss_d / DCAP64LVT
XXFILLER_15_960 vdd_d vss_d / DCAP64LVT
XXFILLER_15_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_18_576 vdd_d vss_d / DCAP64LVT
XXFILLER_15_896 vdd_d vss_d / DCAP64LVT
XXFILLER_15_832 vdd_d vss_d / DCAP64LVT
XXFILLER_15_576 vdd_d vss_d / DCAP64LVT
XXFILLER_15_768 vdd_d vss_d / DCAP64LVT
XXFILLER_15_704 vdd_d vss_d / DCAP64LVT
XXFILLER_15_640 vdd_d vss_d / DCAP64LVT
XXFILLER_17_2216 vdd_d vss_d / DCAP64LVT
XXFILLER_17_2152 vdd_d vss_d / DCAP64LVT
XXFILLER_15_0 vdd_d vss_d / DCAP64LVT
XXFILLER_15_64 vdd_d vss_d / DCAP64LVT
XXFILLER_15_256 vdd_d vss_d / DCAP64LVT
XXFILLER_15_320 vdd_d vss_d / DCAP64LVT
XXFILLER_15_128 vdd_d vss_d / DCAP64LVT
XXFILLER_15_192 vdd_d vss_d / DCAP64LVT
XXFILLER_14_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_14_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_14_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_17_1320 vdd_d vss_d / DCAP64LVT
XXFILLER_17_1256 vdd_d vss_d / DCAP64LVT
XXFILLER_14_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_14_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_14_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_14_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_14_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_14_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_14_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_14_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_14_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_17_384 vdd_d vss_d / DCAP64LVT
XXFILLER_17_448 vdd_d vss_d / DCAP64LVT
XXFILLER_17_320 vdd_d vss_d / DCAP64LVT
XXFILLER_14_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_14_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_14_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_14_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_14_448 vdd_d vss_d / DCAP64LVT
XXFILLER_14_512 vdd_d vss_d / DCAP64LVT
XXFILLER_14_704 vdd_d vss_d / DCAP64LVT
XXFILLER_14_576 vdd_d vss_d / DCAP64LVT
XXFILLER_14_640 vdd_d vss_d / DCAP64LVT
XXFILLER_14_256 vdd_d vss_d / DCAP64LVT
XXFILLER_16_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_14_192 vdd_d vss_d / DCAP64LVT
XXFILLER_14_128 vdd_d vss_d / DCAP64LVT
XXFILLER_13_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_13_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_14_768 vdd_d vss_d / DCAP64LVT
XXFILLER_14_832 vdd_d vss_d / DCAP64LVT
XXFILLER_14_960 vdd_d vss_d / DCAP64LVT
XXFILLER_14_896 vdd_d vss_d / DCAP64LVT
XXFILLER_13_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_13_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_16_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_16_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_13_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_14_64 vdd_d vss_d / DCAP64LVT
XXFILLER_13_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_13_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_13_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_13_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_14_0 vdd_d vss_d / DCAP64LVT
XXFILLER_13_512 vdd_d vss_d / DCAP64LVT
XXFILLER_13_704 vdd_d vss_d / DCAP64LVT
XXFILLER_16_512 vdd_d vss_d / DCAP64LVT
XXFILLER_16_448 vdd_d vss_d / DCAP64LVT
XXFILLER_13_896 vdd_d vss_d / DCAP64LVT
XXFILLER_13_640 vdd_d vss_d / DCAP64LVT
XXFILLER_13_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_13_832 vdd_d vss_d / DCAP64LVT
XXFILLER_13_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_13_960 vdd_d vss_d / DCAP64LVT
XXFILLER_13_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_13_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_13_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_13_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_13_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_13_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_15_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_15_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_13_64 vdd_d vss_d / DCAP64LVT
XXFILLER_13_0 vdd_d vss_d / DCAP64LVT
XXFILLER_13_448 vdd_d vss_d / DCAP64LVT
XXFILLER_13_192 vdd_d vss_d / DCAP64LVT
XXFILLER_13_128 vdd_d vss_d / DCAP64LVT
XXFILLER_13_256 vdd_d vss_d / DCAP64LVT
XXFILLER_13_576 vdd_d vss_d / DCAP64LVT
XXFILLER_13_768 vdd_d vss_d / DCAP64LVT
XXFILLER_15_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_12_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_15_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_12_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_12_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_12_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_12_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_12_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_12_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_12_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_12_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_12_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_15_448 vdd_d vss_d / DCAP64LVT
XXFILLER_12_896 vdd_d vss_d / DCAP64LVT
XXFILLER_15_384 vdd_d vss_d / DCAP64LVT
XXFILLER_12_960 vdd_d vss_d / DCAP64LVT
XXFILLER_12_256 vdd_d vss_d / DCAP64LVT
XXFILLER_12_512 vdd_d vss_d / DCAP64LVT
XXFILLER_12_448 vdd_d vss_d / DCAP64LVT
XXFILLER_12_320 vdd_d vss_d / DCAP64LVT
XXFILLER_12_384 vdd_d vss_d / DCAP64LVT
XXFILLER_12_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_12_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_12_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_12_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_12_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_14_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_12_64 vdd_d vss_d / DCAP64LVT
XXFILLER_14_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_11_1758 vdd_d vss_d / DCAP64LVT
XXFILLER_11_1822 vdd_d vss_d / DCAP64LVT
XXFILLER_12_832 vdd_d vss_d / DCAP64LVT
XXFILLER_11_2014 vdd_d vss_d / DCAP64LVT
XXFILLER_12_576 vdd_d vss_d / DCAP64LVT
XXFILLER_11_1886 vdd_d vss_d / DCAP64LVT
XXFILLER_11_1950 vdd_d vss_d / DCAP64LVT
XXFILLER_12_704 vdd_d vss_d / DCAP64LVT
XXFILLER_12_640 vdd_d vss_d / DCAP64LVT
XXFILLER_12_768 vdd_d vss_d / DCAP64LVT
XXFILLER_11_926 vdd_d vss_d / DCAP64LVT
XXFILLER_11_1054 vdd_d vss_d / DCAP64LVT
XXFILLER_11_990 vdd_d vss_d / DCAP64LVT
XXFILLER_11_1118 vdd_d vss_d / DCAP64LVT
XXFILLER_11_2078 vdd_d vss_d / DCAP64LVT
XXFILLER_11_2270 vdd_d vss_d / DCAP64LVT
XXFILLER_11_2206 vdd_d vss_d / DCAP64LVT
XXFILLER_11_2142 vdd_d vss_d / DCAP64LVT
XXFILLER_11_1566 vdd_d vss_d / DCAP64LVT
XXFILLER_14_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_14_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_11_862 vdd_d vss_d / DCAP64LVT
XXFILLER_12_0 vdd_d vss_d / DCAP64LVT
XXFILLER_14_384 vdd_d vss_d / DCAP64LVT
XXFILLER_11_670 vdd_d vss_d / DCAP64LVT
XXFILLER_14_320 vdd_d vss_d / DCAP64LVT
XXFILLER_11_128 vdd_d vss_d / DCAP64LVT
XXFILLER_11_192 vdd_d vss_d / DCAP64LVT
XXFILLER_11_384 vdd_d vss_d / DCAP64LVT
XXFILLER_11_1182 vdd_d vss_d / DCAP64LVT
XXFILLER_11_256 vdd_d vss_d / DCAP64LVT
XXFILLER_11_320 vdd_d vss_d / DCAP64LVT
XXFILLER_11_1310 vdd_d vss_d / DCAP64LVT
XXFILLER_11_1246 vdd_d vss_d / DCAP64LVT
XXFILLER_11_1374 vdd_d vss_d / DCAP64LVT
XXFILLER_11_1502 vdd_d vss_d / DCAP64LVT
XXFILLER_11_1438 vdd_d vss_d / DCAP64LVT
XXFILLER_13_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_13_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_10_1645 vdd_d vss_d / DCAP64LVT
XXFILLER_10_1773 vdd_d vss_d / DCAP64LVT
XXFILLER_10_1901 vdd_d vss_d / DCAP64LVT
XXFILLER_10_1581 vdd_d vss_d / DCAP64LVT
XXFILLER_10_1709 vdd_d vss_d / DCAP64LVT
XXFILLER_11_448 vdd_d vss_d / DCAP64LVT
XXFILLER_10_1837 vdd_d vss_d / DCAP64LVT
XXFILLER_11_606 vdd_d vss_d / DCAP64LVT
XXFILLER_11_542 vdd_d vss_d / DCAP64LVT
XXFILLER_13_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_10_1057 vdd_d vss_d / DCAP64LVT
XXFILLER_10_993 vdd_d vss_d / DCAP64LVT
XXFILLER_10_1185 vdd_d vss_d / DCAP64LVT
XXFILLER_10_1121 vdd_d vss_d / DCAP64LVT
XXFILLER_10_2285 vdd_d vss_d / DCAP64LVT
XXFILLER_10_2221 vdd_d vss_d / DCAP64LVT
XXFILLER_10_1261 vdd_d vss_d / DCAP64LVT
XXFILLER_10_2029 vdd_d vss_d / DCAP64LVT
XXFILLER_10_1965 vdd_d vss_d / DCAP64LVT
XXFILLER_10_2157 vdd_d vss_d / DCAP64LVT
XXFILLER_10_2093 vdd_d vss_d / DCAP64LVT
XXFILLER_10_192 vdd_d vss_d / DCAP64LVT
XXFILLER_13_384 vdd_d vss_d / DCAP64LVT
XXFILLER_13_320 vdd_d vss_d / DCAP64LVT
XXFILLER_10_128 vdd_d vss_d / DCAP64LVT
XXFILLER_10_64 vdd_d vss_d / DCAP64LVT
XXFILLER_10_320 vdd_d vss_d / DCAP64LVT
XXFILLER_10_256 vdd_d vss_d / DCAP64LVT
XXFILLER_10_929 vdd_d vss_d / DCAP64LVT
XXFILLER_10_1325 vdd_d vss_d / DCAP64LVT
XXFILLER_10_1389 vdd_d vss_d / DCAP64LVT
XXFILLER_10_865 vdd_d vss_d / DCAP64LVT
XXFILLER_9_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_12_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_12_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_10_512 vdd_d vss_d / DCAP64LVT
XXFILLER_10_384 vdd_d vss_d / DCAP64LVT
XXFILLER_10_576 vdd_d vss_d / DCAP64LVT
XXFILLER_10_448 vdd_d vss_d / DCAP64LVT
XXFILLER_10_704 vdd_d vss_d / DCAP64LVT
XXFILLER_10_640 vdd_d vss_d / DCAP64LVT
XXFILLER_12_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_12_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_12_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_9_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_9_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_9_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_9_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_9_832 vdd_d vss_d / DCAP64LVT
XXFILLER_9_896 vdd_d vss_d / DCAP64LVT
XXFILLER_9_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_9_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_9_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_9_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_9_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_12_192 vdd_d vss_d / DCAP64LVT
XXFILLER_12_128 vdd_d vss_d / DCAP64LVT
XXFILLER_9_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_9_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_9_128 vdd_d vss_d / DCAP64LVT
XXFILLER_9_64 vdd_d vss_d / DCAP64LVT
XXFILLER_9_0 vdd_d vss_d / DCAP64LVT
XXFILLER_9_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_9_192 vdd_d vss_d / DCAP64LVT
XXFILLER_9_960 vdd_d vss_d / DCAP64LVT
XXFILLER_9_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_8_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_8_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_8_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_9_256 vdd_d vss_d / DCAP64LVT
XXFILLER_9_320 vdd_d vss_d / DCAP64LVT
XXFILLER_9_448 vdd_d vss_d / DCAP64LVT
XXFILLER_9_384 vdd_d vss_d / DCAP64LVT
XXFILLER_11_1694 vdd_d vss_d / DCAP64LVT
XXFILLER_11_1630 vdd_d vss_d / DCAP64LVT
XXFILLER_8_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_8_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_8_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_9_640 vdd_d vss_d / DCAP64LVT
XXFILLER_9_576 vdd_d vss_d / DCAP64LVT
XXFILLER_9_512 vdd_d vss_d / DCAP64LVT
XXFILLER_11_798 vdd_d vss_d / DCAP64LVT
XXFILLER_11_734 vdd_d vss_d / DCAP64LVT
XXFILLER_8_896 vdd_d vss_d / DCAP64LVT
XXFILLER_8_640 vdd_d vss_d / DCAP64LVT
XXFILLER_8_704 vdd_d vss_d / DCAP64LVT
XXFILLER_8_768 vdd_d vss_d / DCAP64LVT
XXFILLER_8_832 vdd_d vss_d / DCAP64LVT
XXFILLER_8_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_8_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_8_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_8_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_8_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_8_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_11_64 vdd_d vss_d / DCAP64LVT
XXFILLER_11_0 vdd_d vss_d / DCAP64LVT
XXFILLER_8_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_8_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_8_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_8_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_8_960 vdd_d vss_d / DCAP64LVT
XXFILLER_8_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_8_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_8_576 vdd_d vss_d / DCAP64LVT
XXFILLER_8_192 vdd_d vss_d / DCAP64LVT
XXFILLER_8_64 vdd_d vss_d / DCAP64LVT
XXFILLER_8_0 vdd_d vss_d / DCAP64LVT
XXFILLER_8_320 vdd_d vss_d / DCAP64LVT
XXFILLER_8_256 vdd_d vss_d / DCAP64LVT
XXFILLER_8_384 vdd_d vss_d / DCAP64LVT
XXFILLER_7_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_7_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_10_1517 vdd_d vss_d / DCAP64LVT
XXFILLER_10_1453 vdd_d vss_d / DCAP64LVT
XXFILLER_8_128 vdd_d vss_d / DCAP64LVT
XXFILLER_7_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_7_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_7_704 vdd_d vss_d / DCAP64LVT
XXFILLER_7_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_7_640 vdd_d vss_d / DCAP64LVT
XXFILLER_7_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_7_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_7_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_7_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_7_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_7_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_7_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_7_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_7_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_10_0 vdd_d vss_d / DCAP64LVT
XXFILLER_9_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_7_832 vdd_d vss_d / DCAP64LVT
XXFILLER_7_896 vdd_d vss_d / DCAP64LVT
XXFILLER_7_576 vdd_d vss_d / DCAP64LVT
XXFILLER_7_512 vdd_d vss_d / DCAP64LVT
XXFILLER_7_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_7_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_7_960 vdd_d vss_d / DCAP64LVT
XXFILLER_7_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_7_448 vdd_d vss_d / DCAP64LVT
XXFILLER_7_384 vdd_d vss_d / DCAP64LVT
XXFILLER_7_192 vdd_d vss_d / DCAP64LVT
XXFILLER_6_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_6_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_6_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_6_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_7_0 vdd_d vss_d / DCAP64LVT
XXFILLER_9_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_7_128 vdd_d vss_d / DCAP64LVT
XXFILLER_7_64 vdd_d vss_d / DCAP64LVT
XXFILLER_7_768 vdd_d vss_d / DCAP64LVT
XXFILLER_9_768 vdd_d vss_d / DCAP64LVT
XXFILLER_6_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_6_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_9_704 vdd_d vss_d / DCAP64LVT
XXFILLER_6_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_6_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_6_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_6_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_6_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_6_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_6_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_6_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_6_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_6_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_6_896 vdd_d vss_d / DCAP64LVT
XXFILLER_6_832 vdd_d vss_d / DCAP64LVT
XXFILLER_6_512 vdd_d vss_d / DCAP64LVT
XXFILLER_6_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_6_448 vdd_d vss_d / DCAP64LVT
XXFILLER_6_704 vdd_d vss_d / DCAP64LVT
XXFILLER_6_576 vdd_d vss_d / DCAP64LVT
XXFILLER_6_384 vdd_d vss_d / DCAP64LVT
XXFILLER_6_768 vdd_d vss_d / DCAP64LVT
XXFILLER_6_640 vdd_d vss_d / DCAP64LVT
XXFILLER_6_960 vdd_d vss_d / DCAP64LVT
XXFILLER_6_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_8_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_8_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_6_0 vdd_d vss_d / DCAP64LVT
XXFILLER_6_192 vdd_d vss_d / DCAP64LVT
XXFILLER_5_1851 vdd_d vss_d / DCAP64LVT
XXFILLER_5_1915 vdd_d vss_d / DCAP64LVT
XXFILLER_5_1787 vdd_d vss_d / DCAP64LVT
XXFILLER_5_2043 vdd_d vss_d / DCAP64LVT
XXFILLER_5_1979 vdd_d vss_d / DCAP64LVT
XXFILLER_6_320 vdd_d vss_d / DCAP64LVT
XXFILLER_6_256 vdd_d vss_d / DCAP64LVT
XXFILLER_8_512 vdd_d vss_d / DCAP64LVT
XXFILLER_5_1595 vdd_d vss_d / DCAP64LVT
XXFILLER_8_448 vdd_d vss_d / DCAP64LVT
XXFILLER_5_891 vdd_d vss_d / DCAP64LVT
XXFILLER_5_1019 vdd_d vss_d / DCAP64LVT
XXFILLER_5_1147 vdd_d vss_d / DCAP64LVT
XXFILLER_5_955 vdd_d vss_d / DCAP64LVT
XXFILLER_5_2107 vdd_d vss_d / DCAP64LVT
XXFILLER_5_1083 vdd_d vss_d / DCAP64LVT
XXFILLER_5_2171 vdd_d vss_d / DCAP64LVT
XXFILLER_5_2235 vdd_d vss_d / DCAP64LVT
XXFILLER_7_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_5_256 vdd_d vss_d / DCAP64LVT
XXFILLER_5_192 vdd_d vss_d / DCAP64LVT
XXFILLER_5_1531 vdd_d vss_d / DCAP64LVT
XXFILLER_5_1467 vdd_d vss_d / DCAP64LVT
XXFILLER_5_320 vdd_d vss_d / DCAP64LVT
XXFILLER_5_1275 vdd_d vss_d / DCAP64LVT
XXFILLER_5_1211 vdd_d vss_d / DCAP64LVT
XXFILLER_5_1403 vdd_d vss_d / DCAP64LVT
XXFILLER_5_1339 vdd_d vss_d / DCAP64LVT
XXFILLER_5_0 vdd_d vss_d / DCAP64LVT
XXFILLER_5_64 vdd_d vss_d / DCAP64LVT
XXFILLER_5_429 vdd_d vss_d / DCAP64LVT
XXFILLER_5_493 vdd_d vss_d / DCAP64LVT
XXFILLER_7_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_7_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_4_1888 vdd_d vss_d / DCAP64LVT
XXFILLER_4_1824 vdd_d vss_d / DCAP64LVT
XXFILLER_5_621 vdd_d vss_d / DCAP64LVT
XXFILLER_5_557 vdd_d vss_d / DCAP64LVT
XXFILLER_5_685 vdd_d vss_d / DCAP64LVT
XXFILLER_7_320 vdd_d vss_d / DCAP64LVT
XXFILLER_7_256 vdd_d vss_d / DCAP64LVT
XXFILLER_4_928 vdd_d vss_d / DCAP64LVT
XXFILLER_4_1632 vdd_d vss_d / DCAP64LVT
XXFILLER_4_1696 vdd_d vss_d / DCAP64LVT
XXFILLER_4_1568 vdd_d vss_d / DCAP64LVT
XXFILLER_4_2080 vdd_d vss_d / DCAP64LVT
XXFILLER_4_2144 vdd_d vss_d / DCAP64LVT
XXFILLER_4_1952 vdd_d vss_d / DCAP64LVT
XXFILLER_4_2016 vdd_d vss_d / DCAP64LVT
XXFILLER_4_2272 vdd_d vss_d / DCAP64LVT
XXFILLER_4_2208 vdd_d vss_d / DCAP64LVT
XXFILLER_4_992 vdd_d vss_d / DCAP64LVT
XXFILLER_4_1184 vdd_d vss_d / DCAP64LVT
XXFILLER_4_1056 vdd_d vss_d / DCAP64LVT
XXFILLER_4_1120 vdd_d vss_d / DCAP64LVT
XXFILLER_4_1312 vdd_d vss_d / DCAP64LVT
XXFILLER_4_1440 vdd_d vss_d / DCAP64LVT
XXFILLER_4_1376 vdd_d vss_d / DCAP64LVT
XXFILLER_4_1248 vdd_d vss_d / DCAP64LVT
XXFILLER_4_320 vdd_d vss_d / DCAP64LVT
XXFILLER_6_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_4_256 vdd_d vss_d / DCAP64LVT
XXFILLER_4_1504 vdd_d vss_d / DCAP64LVT
XXFILLER_6_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_3_2148 vdd_d vss_d / DCAP64LVT
XXFILLER_3_1892 vdd_d vss_d / DCAP64LVT
XXFILLER_3_2020 vdd_d vss_d / DCAP64LVT
XXFILLER_3_1956 vdd_d vss_d / DCAP64LVT
XXFILLER_3_2084 vdd_d vss_d / DCAP64LVT
XXFILLER_4_672 vdd_d vss_d / DCAP64LVT
XXFILLER_4_416 vdd_d vss_d / DCAP64LVT
XXFILLER_4_480 vdd_d vss_d / DCAP64LVT
XXFILLER_4_544 vdd_d vss_d / DCAP64LVT
XXFILLER_4_608 vdd_d vss_d / DCAP64LVT
XXFILLER_4_736 vdd_d vss_d / DCAP64LVT
XXFILLER_6_128 vdd_d vss_d / DCAP64LVT
XXFILLER_3_996 vdd_d vss_d / DCAP64LVT
XXFILLER_6_64 vdd_d vss_d / DCAP64LVT
XXFILLER_3_1060 vdd_d vss_d / DCAP64LVT
XXFILLER_3_1124 vdd_d vss_d / DCAP64LVT
XXFILLER_4_64 vdd_d vss_d / DCAP64LVT
XXFILLER_4_0 vdd_d vss_d / DCAP64LVT
XXFILLER_3_2212 vdd_d vss_d / DCAP64LVT
XXFILLER_3_2276 vdd_d vss_d / DCAP64LVT
XXFILLER_3_1252 vdd_d vss_d / DCAP64LVT
XXFILLER_3_1188 vdd_d vss_d / DCAP64LVT
XXFILLER_5_1723 vdd_d vss_d / DCAP64LVT
XXFILLER_5_1659 vdd_d vss_d / DCAP64LVT
XXFILLER_3_1700 vdd_d vss_d / DCAP64LVT
XXFILLER_3_1508 vdd_d vss_d / DCAP64LVT
XXFILLER_3_1316 vdd_d vss_d / DCAP64LVT
XXFILLER_3_1444 vdd_d vss_d / DCAP64LVT
XXFILLER_3_1636 vdd_d vss_d / DCAP64LVT
XXFILLER_3_1380 vdd_d vss_d / DCAP64LVT
XXFILLER_3_1572 vdd_d vss_d / DCAP64LVT
XXFILLER_5_827 vdd_d vss_d / DCAP64LVT
XXFILLER_2_1954 vdd_d vss_d / DCAP64LVT
XXFILLER_5_763 vdd_d vss_d / DCAP64LVT
XXFILLER_2_2018 vdd_d vss_d / DCAP64LVT
XXFILLER_2_2146 vdd_d vss_d / DCAP64LVT
XXFILLER_3_548 vdd_d vss_d / DCAP64LVT
XXFILLER_2_2082 vdd_d vss_d / DCAP64LVT
XXFILLER_3_484 vdd_d vss_d / DCAP64LVT
XXFILLER_3_740 vdd_d vss_d / DCAP64LVT
XXFILLER_3_612 vdd_d vss_d / DCAP64LVT
XXFILLER_3_420 vdd_d vss_d / DCAP64LVT
XXFILLER_3_804 vdd_d vss_d / DCAP64LVT
XXFILLER_3_676 vdd_d vss_d / DCAP64LVT
XXFILLER_3_320 vdd_d vss_d / DCAP64LVT
XXFILLER_5_128 vdd_d vss_d / DCAP64LVT
XXFILLER_2_1058 vdd_d vss_d / DCAP64LVT
XXFILLER_2_994 vdd_d vss_d / DCAP64LVT
XXFILLER_2_1122 vdd_d vss_d / DCAP64LVT
XXFILLER_2_1250 vdd_d vss_d / DCAP64LVT
XXFILLER_2_1186 vdd_d vss_d / DCAP64LVT
XXFILLER_2_1890 vdd_d vss_d / DCAP64LVT
XXFILLER_3_64 vdd_d vss_d / DCAP64LVT
XXFILLER_3_0 vdd_d vss_d / DCAP64LVT
XXFILLER_2_2210 vdd_d vss_d / DCAP64LVT
XXFILLER_2_2274 vdd_d vss_d / DCAP64LVT
XXFILLER_3_128 vdd_d vss_d / DCAP64LVT
XXFILLER_2_1634 vdd_d vss_d / DCAP64LVT
XXFILLER_4_1760 vdd_d vss_d / DCAP64LVT
XXFILLER_2_1442 vdd_d vss_d / DCAP64LVT
XXFILLER_2_1506 vdd_d vss_d / DCAP64LVT
XXFILLER_2_1314 vdd_d vss_d / DCAP64LVT
XXFILLER_2_1378 vdd_d vss_d / DCAP64LVT
XXFILLER_2_1698 vdd_d vss_d / DCAP64LVT
XXFILLER_2_1570 vdd_d vss_d / DCAP64LVT
XXFILLER_4_864 vdd_d vss_d / DCAP64LVT
XXFILLER_4_800 vdd_d vss_d / DCAP64LVT
XXFILLER_4_192 vdd_d vss_d / DCAP64LVT
XXFILLER_4_128 vdd_d vss_d / DCAP64LVT
XXFILLER_1_2239 vdd_d vss_d / DCAP64LVT
XXFILLER_1_2175 vdd_d vss_d / DCAP64LVT
XXFILLER_2_543 vdd_d vss_d / DCAP64LVT
XXFILLER_2_384 vdd_d vss_d / DCAP64LVT
XXFILLER_3_1828 vdd_d vss_d / DCAP64LVT
XXFILLER_1_1215 vdd_d vss_d / DCAP64LVT
XXFILLER_3_1764 vdd_d vss_d / DCAP64LVT
XXFILLER_1_1279 vdd_d vss_d / DCAP64LVT
XXFILLER_1_1407 vdd_d vss_d / DCAP64LVT
XXFILLER_1_1343 vdd_d vss_d / DCAP64LVT
XXFILLER_2_0 vdd_d vss_d / DCAP64LVT
XXFILLER_2_64 vdd_d vss_d / DCAP64LVT
XXFILLER_2_192 vdd_d vss_d / DCAP64LVT
XXFILLER_2_128 vdd_d vss_d / DCAP64LVT
XXFILLER_1_2047 vdd_d vss_d / DCAP64LVT
XXFILLER_1_2111 vdd_d vss_d / DCAP64LVT
XXFILLER_3_932 vdd_d vss_d / DCAP64LVT
XXFILLER_1_512 vdd_d vss_d / DCAP64LVT
XXFILLER_3_868 vdd_d vss_d / DCAP64LVT
XXFILLER_1_576 vdd_d vss_d / DCAP64LVT
XXFILLER_1_704 vdd_d vss_d / DCAP64LVT
XXFILLER_1_1599 vdd_d vss_d / DCAP64LVT
XXFILLER_1_640 vdd_d vss_d / DCAP64LVT
XXFILLER_1_1535 vdd_d vss_d / DCAP64LVT
XXFILLER_1_1791 vdd_d vss_d / DCAP64LVT
XXFILLER_1_1663 vdd_d vss_d / DCAP64LVT
XXFILLER_1_1471 vdd_d vss_d / DCAP64LVT
XXFILLER_1_1855 vdd_d vss_d / DCAP64LVT
XXFILLER_1_1727 vdd_d vss_d / DCAP64LVT
XXFILLER_1_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_3_256 vdd_d vss_d / DCAP64LVT
XXFILLER_0_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_3_192 vdd_d vss_d / DCAP64LVT
XXFILLER_0_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_0_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_1_448 vdd_d vss_d / DCAP64LVT
XXFILLER_1_895 vdd_d vss_d / DCAP64LVT
XXFILLER_1_831 vdd_d vss_d / DCAP64LVT
XXFILLER_1_320 vdd_d vss_d / DCAP64LVT
XXFILLER_1_959 vdd_d vss_d / DCAP64LVT
XXFILLER_1_384 vdd_d vss_d / DCAP64LVT
XXFILLER_2_1826 vdd_d vss_d / DCAP64LVT
XXFILLER_0_640 vdd_d vss_d / DCAP64LVT
XXFILLER_2_1762 vdd_d vss_d / DCAP64LVT
XXFILLER_0_576 vdd_d vss_d / DCAP64LVT
XXFILLER_0_704 vdd_d vss_d / DCAP64LVT
XXFILLER_0_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_0_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_0_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_0_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_0_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_0_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_0_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_0_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_0_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_0_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_2_930 vdd_d vss_d / DCAP64LVT
XXFILLER_2_866 vdd_d vss_d / DCAP64LVT
XXFILLER_0_896 vdd_d vss_d / DCAP64LVT
XXFILLER_0_384 vdd_d vss_d / DCAP64LVT
XXFILLER_0_832 vdd_d vss_d / DCAP64LVT
XXFILLER_0_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_0_960 vdd_d vss_d / DCAP64LVT
XXFILLER_0_768 vdd_d vss_d / DCAP64LVT
XXFILLER_0_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_0_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_0_512 vdd_d vss_d / DCAP64LVT
XXFILLER_0_448 vdd_d vss_d / DCAP64LVT
XXFILLER_2_626 vdd_d vss_d / DCAP64LVT
XXFILLER_0_128 vdd_d vss_d / DCAP64LVT
XXFILLER_0_64 vdd_d vss_d / DCAP64LVT
XXFILLER_0_0 vdd_d vss_d / DCAP64LVT
XXFILLER_0_192 vdd_d vss_d / DCAP64LVT
XXFILLER_2_320 vdd_d vss_d / DCAP64LVT
XXFILLER_2_256 vdd_d vss_d / DCAP64LVT
XXFILLER_1_1983 vdd_d vss_d / DCAP64LVT
XXFILLER_1_1919 vdd_d vss_d / DCAP64LVT
XXFILLER_1_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_1_1023 vdd_d vss_d / DCAP64LVT
XXFILLER_1_192 vdd_d vss_d / DCAP64LVT
XXFILLER_1_128 vdd_d vss_d / DCAP64LVT
XXFILLER_1_64 vdd_d vss_d / DCAP64LVT
XXFILLER_1_0 vdd_d vss_d / DCAP64LVT
XXFILLER_1_256 vdd_d vss_d / DCAP64LVT
XXFILLER_0_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_0_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_0_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_0_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_0_320 vdd_d vss_d / DCAP64LVT
XXFILLER_0_256 vdd_d vss_d / DCAP64LVT
XXFILLER_17_192 vdd_d vss_d / DCAP64LVT
XXFILLER_9_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_9_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_17_64 vdd_d vss_d / DCAP64LVT
XXFILLER_17_0 vdd_d vss_d / DCAP64LVT
XXFILLER_9_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_9_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_17_256 vdd_d vss_d / DCAP64LVT
XXFILLER_17_128 vdd_d vss_d / DCAP64LVT
XXFILLER_20_1039 vdd_d vss_d / DCAP64LVT
XXFILLER_20_960 vdd_d vss_d / DCAP64LVT
XXFILLER_20_896 vdd_d vss_d / DCAP64LVT
XXFILLER_20_832 vdd_d vss_d / DCAP64LVT
XXFILLER_20_768 vdd_d vss_d / DCAP64LVT
XXFILLER_20_704 vdd_d vss_d / DCAP64LVT
XXFILLER_20_640 vdd_d vss_d / DCAP64LVT
XXFILLER_20_576 vdd_d vss_d / DCAP64LVT
XXFILLER_20_512 vdd_d vss_d / DCAP64LVT
XXFILLER_20_448 vdd_d vss_d / DCAP64LVT
XXFILLER_20_384 vdd_d vss_d / DCAP64LVT
XXFILLER_20_192 vdd_d vss_d / DCAP64LVT
XXFILLER_20_128 vdd_d vss_d / DCAP64LVT
XXFILLER_17_936 vdd_d vss_d / DCAP64LVT
XXFILLER_17_872 vdd_d vss_d / DCAP64LVT
XXFILLER_17_1000 vdd_d vss_d / DCAP64LVT
XXFILLER_17_1064 vdd_d vss_d / DCAP64LVT
XXFILLER_17_1192 vdd_d vss_d / DCAP64LVT
XXFILLER_17_1128 vdd_d vss_d / DCAP64LVT
XXFILLER_17_552 vdd_d vss_d / DCAP64LVT
XXFILLER_17_680 vdd_d vss_d / DCAP64LVT
XXFILLER_17_616 vdd_d vss_d / DCAP64LVT
XXFILLER_17_744 vdd_d vss_d / DCAP64LVT
XXFILLER_17_1704 vdd_d vss_d / DCAP64LVT
XXFILLER_17_1832 vdd_d vss_d / DCAP64LVT
XXFILLER_17_1768 vdd_d vss_d / DCAP64LVT
XXFILLER_17_1896 vdd_d vss_d / DCAP64LVT
XXFILLER_17_2024 vdd_d vss_d / DCAP64LVT
XXFILLER_17_1960 vdd_d vss_d / DCAP64LVT
XXFILLER_17_2088 vdd_d vss_d / DCAP64LVT
XXFILLER_17_1384 vdd_d vss_d / DCAP64LVT
XXFILLER_17_1448 vdd_d vss_d / DCAP64LVT
XXFILLER_17_1576 vdd_d vss_d / DCAP64LVT
XXFILLER_17_1512 vdd_d vss_d / DCAP64LVT
XXFILLER_17_1640 vdd_d vss_d / DCAP64LVT
XXFILLER_18_0 vdd_d vss_d / DCAP64LVT
XXFILLER_18_128 vdd_d vss_d / DCAP64LVT
XXFILLER_18_64 vdd_d vss_d / DCAP64LVT
XXFILLER_18_192 vdd_d vss_d / DCAP64LVT
XXFILLER_18_256 vdd_d vss_d / DCAP64LVT
XXFILLER_17_2280 vdd_d vss_d / DCAP64LVT
XXFILLER_18_448 vdd_d vss_d / DCAP64LVT
XXFILLER_18_384 vdd_d vss_d / DCAP64LVT
XXFILLER_18_320 vdd_d vss_d / DCAP64LVT
XXFILLER_18_512 vdd_d vss_d / DCAP64LVT
XXFILLER_18_640 vdd_d vss_d / DCAP64LVT
XXFILLER_18_704 vdd_d vss_d / DCAP64LVT
XXFILLER_18_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_18_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_18_896 vdd_d vss_d / DCAP64LVT
XXFILLER_18_960 vdd_d vss_d / DCAP64LVT
XXFILLER_18_768 vdd_d vss_d / DCAP64LVT
XXFILLER_18_832 vdd_d vss_d / DCAP64LVT
XXFILLER_18_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_18_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_18_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_18_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_18_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_18_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_18_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_18_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_18_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_18_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_18_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_18_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_18_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_18_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_18_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_18_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_18_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_19_192 vdd_d vss_d / DCAP64LVT
XXFILLER_19_256 vdd_d vss_d / DCAP64LVT
XXFILLER_19_64 vdd_d vss_d / DCAP64LVT
XXFILLER_19_128 vdd_d vss_d / DCAP64LVT
XXFILLER_19_384 vdd_d vss_d / DCAP64LVT
XXFILLER_19_320 vdd_d vss_d / DCAP64LVT
XXFILLER_19_448 vdd_d vss_d / DCAP64LVT
XXFILLER_19_0 vdd_d vss_d / DCAP64LVT
XXFILLER_19_994 vdd_d vss_d / DCAP64LVT
XXFILLER_19_1058 vdd_d vss_d / DCAP64LVT
XXFILLER_19_866 vdd_d vss_d / DCAP64LVT
XXFILLER_19_930 vdd_d vss_d / DCAP64LVT
XXFILLER_19_546 vdd_d vss_d / DCAP64LVT
XXFILLER_19_610 vdd_d vss_d / DCAP64LVT
XXFILLER_19_738 vdd_d vss_d / DCAP64LVT
XXFILLER_19_674 vdd_d vss_d / DCAP64LVT
XXFILLER_19_802 vdd_d vss_d / DCAP64LVT
XXFILLER_19_1683 vdd_d vss_d / DCAP64LVT
XXFILLER_19_1747 vdd_d vss_d / DCAP64LVT
XXFILLER_19_1619 vdd_d vss_d / DCAP64LVT
XXFILLER_19_1875 vdd_d vss_d / DCAP64LVT
XXFILLER_19_1811 vdd_d vss_d / DCAP64LVT
XXFILLER_19_1939 vdd_d vss_d / DCAP64LVT
XXFILLER_19_2003 vdd_d vss_d / DCAP64LVT
XXFILLER_19_2131 vdd_d vss_d / DCAP64LVT
XXFILLER_19_2067 vdd_d vss_d / DCAP64LVT
XXFILLER_19_2195 vdd_d vss_d / DCAP64LVT
XXFILLER_19_2259 vdd_d vss_d / DCAP64LVT
XXFILLER_19_1363 vdd_d vss_d / DCAP64LVT
XXFILLER_19_1171 vdd_d vss_d / DCAP64LVT
XXFILLER_19_1235 vdd_d vss_d / DCAP64LVT
XXFILLER_20_1252 vdd_d vss_d / DCAP64LVT
XXFILLER_20_1316 vdd_d vss_d / DCAP64LVT
XXFILLER_20_1380 vdd_d vss_d / DCAP64LVT
XXFILLER_20_1444 vdd_d vss_d / DCAP64LVT
XXFILLER_20_1508 vdd_d vss_d / DCAP64LVT
XXFILLER_20_1621 vdd_d vss_d / DCAP64LVT
XXFILLER_20_1762 vdd_d vss_d / DCAP64LVT
XXFILLER_20_1826 vdd_d vss_d / DCAP64LVT
XXFILLER_20_1890 vdd_d vss_d / DCAP64LVT
XXFILLER_20_1954 vdd_d vss_d / DCAP64LVT
XXFILLER_20_2018 vdd_d vss_d / DCAP64LVT
XXFILLER_20_2082 vdd_d vss_d / DCAP64LVT
XXFILLER_20_2146 vdd_d vss_d / DCAP64LVT
XXFILLER_20_2210 vdd_d vss_d / DCAP64LVT
XXFILLER_20_2274 vdd_d vss_d / DCAP64LVT
XXFILLER_21_0 vdd_d vss_d / DCAP64LVT
XXFILLER_21_64 vdd_d vss_d / DCAP64LVT
XXFILLER_21_128 vdd_d vss_d / DCAP64LVT
XXFILLER_21_192 vdd_d vss_d / DCAP64LVT
XXFILLER_21_256 vdd_d vss_d / DCAP64LVT
XXFILLER_21_320 vdd_d vss_d / DCAP64LVT
XXFILLER_21_384 vdd_d vss_d / DCAP64LVT
XXFILLER_21_470 vdd_d vss_d / DCAP64LVT
XXFILLER_21_534 vdd_d vss_d / DCAP64LVT
XXFILLER_21_598 vdd_d vss_d / DCAP64LVT
XXFILLER_21_662 vdd_d vss_d / DCAP64LVT
XXFILLER_21_726 vdd_d vss_d / DCAP64LVT
XXFILLER_21_790 vdd_d vss_d / DCAP64LVT
XXFILLER_21_854 vdd_d vss_d / DCAP64LVT
XXFILLER_21_918 vdd_d vss_d / DCAP64LVT
XXFILLER_21_982 vdd_d vss_d / DCAP64LVT
XXFILLER_21_1046 vdd_d vss_d / DCAP64LVT
XXFILLER_21_1293 vdd_d vss_d / DCAP64LVT
XXFILLER_21_1357 vdd_d vss_d / DCAP64LVT
XXFILLER_21_1421 vdd_d vss_d / DCAP64LVT
XXFILLER_21_1485 vdd_d vss_d / DCAP64LVT
XXFILLER_21_1614 vdd_d vss_d / DCAP64LVT
XXFILLER_21_1678 vdd_d vss_d / DCAP64LVT
XXFILLER_21_1742 vdd_d vss_d / DCAP64LVT
XXFILLER_21_1806 vdd_d vss_d / DCAP64LVT
XXFILLER_21_1870 vdd_d vss_d / DCAP64LVT
XXFILLER_21_1934 vdd_d vss_d / DCAP64LVT
XXFILLER_21_1998 vdd_d vss_d / DCAP64LVT
XXFILLER_21_2062 vdd_d vss_d / DCAP64LVT
XXFILLER_21_2126 vdd_d vss_d / DCAP64LVT
XXFILLER_21_2190 vdd_d vss_d / DCAP64LVT
XXFILLER_21_2254 vdd_d vss_d / DCAP64LVT
XXFILLER_22_0 vdd_d vss_d / DCAP64LVT
XXFILLER_22_64 vdd_d vss_d / DCAP64LVT
XXFILLER_22_128 vdd_d vss_d / DCAP64LVT
XXFILLER_22_192 vdd_d vss_d / DCAP64LVT
XXFILLER_22_256 vdd_d vss_d / DCAP64LVT
XXFILLER_22_320 vdd_d vss_d / DCAP64LVT
XXFILLER_22_384 vdd_d vss_d / DCAP64LVT
XXFILLER_22_448 vdd_d vss_d / DCAP64LVT
XXFILLER_22_512 vdd_d vss_d / DCAP64LVT
XXFILLER_22_576 vdd_d vss_d / DCAP64LVT
XXFILLER_22_640 vdd_d vss_d / DCAP64LVT
XXFILLER_22_704 vdd_d vss_d / DCAP64LVT
XXFILLER_22_768 vdd_d vss_d / DCAP64LVT
XXFILLER_22_832 vdd_d vss_d / DCAP64LVT
XXFILLER_22_896 vdd_d vss_d / DCAP64LVT
XXFILLER_22_960 vdd_d vss_d / DCAP64LVT
XXFILLER_22_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_22_1160 vdd_d vss_d / DCAP64LVT
XXFILLER_22_1246 vdd_d vss_d / DCAP64LVT
XXFILLER_22_1335 vdd_d vss_d / DCAP64LVT
XXFILLER_22_1399 vdd_d vss_d / DCAP64LVT
XXFILLER_22_1463 vdd_d vss_d / DCAP64LVT
XXFILLER_22_1527 vdd_d vss_d / DCAP64LVT
XXFILLER_22_1591 vdd_d vss_d / DCAP64LVT
XXFILLER_22_1655 vdd_d vss_d / DCAP64LVT
XXFILLER_22_1719 vdd_d vss_d / DCAP64LVT
XXFILLER_22_1783 vdd_d vss_d / DCAP64LVT
XXFILLER_22_1847 vdd_d vss_d / DCAP64LVT
XXFILLER_22_1911 vdd_d vss_d / DCAP64LVT
XXFILLER_22_1975 vdd_d vss_d / DCAP64LVT
XXFILLER_22_2039 vdd_d vss_d / DCAP64LVT
XXFILLER_22_2103 vdd_d vss_d / DCAP64LVT
XXFILLER_22_2167 vdd_d vss_d / DCAP64LVT
XXFILLER_22_2231 vdd_d vss_d / DCAP64LVT
XXFILLER_23_0 vdd_d vss_d / DCAP64LVT
XXFILLER_23_64 vdd_d vss_d / DCAP64LVT
XXFILLER_23_128 vdd_d vss_d / DCAP64LVT
XXFILLER_23_192 vdd_d vss_d / DCAP64LVT
XXFILLER_23_256 vdd_d vss_d / DCAP64LVT
XXFILLER_23_320 vdd_d vss_d / DCAP64LVT
XXFILLER_23_461 vdd_d vss_d / DCAP64LVT
XXFILLER_23_525 vdd_d vss_d / DCAP64LVT
XXFILLER_23_589 vdd_d vss_d / DCAP64LVT
XXFILLER_23_653 vdd_d vss_d / DCAP64LVT
XXFILLER_23_717 vdd_d vss_d / DCAP64LVT
XXFILLER_23_781 vdd_d vss_d / DCAP64LVT
XXFILLER_23_845 vdd_d vss_d / DCAP64LVT
XXFILLER_23_909 vdd_d vss_d / DCAP64LVT
XXFILLER_23_973 vdd_d vss_d / DCAP64LVT
XXFILLER_23_1251 vdd_d vss_d / DCAP64LVT
XXFILLER_23_1364 vdd_d vss_d / DCAP64LVT
XXFILLER_23_1428 vdd_d vss_d / DCAP64LVT
XXFILLER_23_1492 vdd_d vss_d / DCAP64LVT
XXFILLER_23_1556 vdd_d vss_d / DCAP64LVT
XXFILLER_23_1620 vdd_d vss_d / DCAP64LVT
XXFILLER_23_1684 vdd_d vss_d / DCAP64LVT
XXFILLER_23_1777 vdd_d vss_d / DCAP64LVT
XXFILLER_23_1841 vdd_d vss_d / DCAP64LVT
XXFILLER_23_1905 vdd_d vss_d / DCAP64LVT
XXFILLER_23_1969 vdd_d vss_d / DCAP64LVT
XXFILLER_23_2033 vdd_d vss_d / DCAP64LVT
XXFILLER_23_2097 vdd_d vss_d / DCAP64LVT
XXFILLER_23_2161 vdd_d vss_d / DCAP64LVT
XXFILLER_23_2225 vdd_d vss_d / DCAP64LVT
XXFILLER_24_0 vdd_d vss_d / DCAP64LVT
XXFILLER_24_64 vdd_d vss_d / DCAP64LVT
XXFILLER_24_128 vdd_d vss_d / DCAP64LVT
XXFILLER_24_192 vdd_d vss_d / DCAP64LVT
XXFILLER_24_256 vdd_d vss_d / DCAP64LVT
XXFILLER_24_320 vdd_d vss_d / DCAP64LVT
XXFILLER_24_459 vdd_d vss_d / DCAP64LVT
XXFILLER_24_523 vdd_d vss_d / DCAP64LVT
XXFILLER_24_587 vdd_d vss_d / DCAP64LVT
XXFILLER_24_651 vdd_d vss_d / DCAP64LVT
XXFILLER_24_715 vdd_d vss_d / DCAP64LVT
XXFILLER_24_779 vdd_d vss_d / DCAP64LVT
XXFILLER_24_843 vdd_d vss_d / DCAP64LVT
XXFILLER_24_907 vdd_d vss_d / DCAP64LVT
XXFILLER_24_971 vdd_d vss_d / DCAP64LVT
XXFILLER_24_1082 vdd_d vss_d / DCAP64LVT
XXFILLER_24_1146 vdd_d vss_d / DCAP64LVT
XXFILLER_24_1236 vdd_d vss_d / DCAP64LVT
XXFILLER_24_1300 vdd_d vss_d / DCAP64LVT
XXFILLER_24_1364 vdd_d vss_d / DCAP64LVT
XXFILLER_24_1428 vdd_d vss_d / DCAP64LVT
XXFILLER_24_1492 vdd_d vss_d / DCAP64LVT
XXFILLER_24_1556 vdd_d vss_d / DCAP64LVT
XXFILLER_24_1669 vdd_d vss_d / DCAP64LVT
XXFILLER_24_1733 vdd_d vss_d / DCAP64LVT
XXFILLER_24_1797 vdd_d vss_d / DCAP64LVT
XXFILLER_24_1861 vdd_d vss_d / DCAP64LVT
XXFILLER_24_1925 vdd_d vss_d / DCAP64LVT
XXFILLER_24_1989 vdd_d vss_d / DCAP64LVT
XXFILLER_24_2053 vdd_d vss_d / DCAP64LVT
XXFILLER_24_2117 vdd_d vss_d / DCAP64LVT
XXFILLER_24_2181 vdd_d vss_d / DCAP64LVT
XXFILLER_24_2245 vdd_d vss_d / DCAP64LVT
XXFILLER_25_0 vdd_d vss_d / DCAP64LVT
XXFILLER_25_64 vdd_d vss_d / DCAP64LVT
XXFILLER_25_128 vdd_d vss_d / DCAP64LVT
XXFILLER_25_192 vdd_d vss_d / DCAP64LVT
XXFILLER_25_256 vdd_d vss_d / DCAP64LVT
XXFILLER_25_320 vdd_d vss_d / DCAP64LVT
XXFILLER_25_384 vdd_d vss_d / DCAP64LVT
XXFILLER_25_448 vdd_d vss_d / DCAP64LVT
XXFILLER_25_528 vdd_d vss_d / DCAP64LVT
XXFILLER_25_592 vdd_d vss_d / DCAP64LVT
XXFILLER_25_656 vdd_d vss_d / DCAP64LVT
XXFILLER_25_720 vdd_d vss_d / DCAP64LVT
XXFILLER_25_784 vdd_d vss_d / DCAP64LVT
XXFILLER_25_848 vdd_d vss_d / DCAP64LVT
XXFILLER_25_912 vdd_d vss_d / DCAP64LVT
XXFILLER_25_976 vdd_d vss_d / DCAP64LVT
XXFILLER_25_1290 vdd_d vss_d / DCAP64LVT
XXFILLER_25_1354 vdd_d vss_d / DCAP64LVT
XXFILLER_25_1418 vdd_d vss_d / DCAP64LVT
XXFILLER_25_1482 vdd_d vss_d / DCAP64LVT
XXFILLER_25_1546 vdd_d vss_d / DCAP64LVT
XXFILLER_25_1610 vdd_d vss_d / DCAP64LVT
XXFILLER_25_1674 vdd_d vss_d / DCAP64LVT
XXFILLER_25_1738 vdd_d vss_d / DCAP64LVT
XXFILLER_25_1802 vdd_d vss_d / DCAP64LVT
XXFILLER_25_1866 vdd_d vss_d / DCAP64LVT
XXFILLER_25_1930 vdd_d vss_d / DCAP64LVT
XXFILLER_25_1994 vdd_d vss_d / DCAP64LVT
XXFILLER_25_2058 vdd_d vss_d / DCAP64LVT
XXFILLER_25_2122 vdd_d vss_d / DCAP64LVT
XXFILLER_25_2186 vdd_d vss_d / DCAP64LVT
XXFILLER_25_2250 vdd_d vss_d / DCAP64LVT
XXFILLER_26_0 vdd_d vss_d / DCAP64LVT
XXFILLER_26_64 vdd_d vss_d / DCAP64LVT
XXFILLER_26_128 vdd_d vss_d / DCAP64LVT
XXFILLER_26_192 vdd_d vss_d / DCAP64LVT
XXFILLER_26_256 vdd_d vss_d / DCAP64LVT
XXFILLER_26_320 vdd_d vss_d / DCAP64LVT
XXFILLER_26_459 vdd_d vss_d / DCAP64LVT
XXFILLER_26_523 vdd_d vss_d / DCAP64LVT
XXFILLER_26_587 vdd_d vss_d / DCAP64LVT
XXFILLER_26_651 vdd_d vss_d / DCAP64LVT
XXFILLER_26_715 vdd_d vss_d / DCAP64LVT
XXFILLER_26_779 vdd_d vss_d / DCAP64LVT
XXFILLER_26_843 vdd_d vss_d / DCAP64LVT
XXFILLER_26_907 vdd_d vss_d / DCAP64LVT
XXFILLER_26_971 vdd_d vss_d / DCAP64LVT
XXFILLER_26_1089 vdd_d vss_d / DCAP64LVT
XXFILLER_26_1153 vdd_d vss_d / DCAP64LVT
XXFILLER_26_1246 vdd_d vss_d / DCAP64LVT
XXFILLER_26_1310 vdd_d vss_d / DCAP64LVT
XXFILLER_26_1435 vdd_d vss_d / DCAP64LVT
XXFILLER_26_1499 vdd_d vss_d / DCAP64LVT
XXFILLER_26_1563 vdd_d vss_d / DCAP64LVT
XXFILLER_26_1627 vdd_d vss_d / DCAP64LVT
XXFILLER_26_1741 vdd_d vss_d / DCAP64LVT
XXFILLER_26_1805 vdd_d vss_d / DCAP64LVT
XXFILLER_26_1869 vdd_d vss_d / DCAP64LVT
XXFILLER_26_1933 vdd_d vss_d / DCAP64LVT
XXFILLER_26_1997 vdd_d vss_d / DCAP64LVT
XXFILLER_26_2061 vdd_d vss_d / DCAP64LVT
XXFILLER_26_2125 vdd_d vss_d / DCAP64LVT
XXFILLER_26_2189 vdd_d vss_d / DCAP64LVT
XXFILLER_26_2253 vdd_d vss_d / DCAP64LVT
XXFILLER_27_0 vdd_d vss_d / DCAP64LVT
XXFILLER_27_64 vdd_d vss_d / DCAP64LVT
XXFILLER_27_128 vdd_d vss_d / DCAP64LVT
XXFILLER_27_192 vdd_d vss_d / DCAP64LVT
XXFILLER_27_256 vdd_d vss_d / DCAP64LVT
XXFILLER_27_320 vdd_d vss_d / DCAP64LVT
XXFILLER_27_504 vdd_d vss_d / DCAP64LVT
XXFILLER_27_568 vdd_d vss_d / DCAP64LVT
XXFILLER_27_632 vdd_d vss_d / DCAP64LVT
XXFILLER_27_696 vdd_d vss_d / DCAP64LVT
XXFILLER_27_760 vdd_d vss_d / DCAP64LVT
XXFILLER_27_824 vdd_d vss_d / DCAP64LVT
XXFILLER_27_888 vdd_d vss_d / DCAP64LVT
XXFILLER_27_1074 vdd_d vss_d / DCAP64LVT
XXFILLER_27_1138 vdd_d vss_d / DCAP64LVT
XXFILLER_27_1202 vdd_d vss_d / DCAP64LVT
XXFILLER_27_1266 vdd_d vss_d / DCAP64LVT
XXFILLER_27_1330 vdd_d vss_d / DCAP64LVT
XXFILLER_27_1394 vdd_d vss_d / DCAP64LVT
XXFILLER_27_1458 vdd_d vss_d / DCAP64LVT
XXFILLER_27_1522 vdd_d vss_d / DCAP64LVT
XXFILLER_27_1586 vdd_d vss_d / DCAP64LVT
XXFILLER_27_1650 vdd_d vss_d / DCAP64LVT
XXFILLER_27_1714 vdd_d vss_d / DCAP64LVT
XXFILLER_27_1840 vdd_d vss_d / DCAP64LVT
XXFILLER_27_1904 vdd_d vss_d / DCAP64LVT
XXFILLER_27_1968 vdd_d vss_d / DCAP64LVT
XXFILLER_27_2032 vdd_d vss_d / DCAP64LVT
XXFILLER_27_2096 vdd_d vss_d / DCAP64LVT
XXFILLER_27_2160 vdd_d vss_d / DCAP64LVT
XXFILLER_27_2224 vdd_d vss_d / DCAP64LVT
XXFILLER_28_0 vdd_d vss_d / DCAP64LVT
XXFILLER_28_64 vdd_d vss_d / DCAP64LVT
XXFILLER_28_128 vdd_d vss_d / DCAP64LVT
XXFILLER_28_192 vdd_d vss_d / DCAP64LVT
XXFILLER_28_256 vdd_d vss_d / DCAP64LVT
XXFILLER_28_320 vdd_d vss_d / DCAP64LVT
XXFILLER_28_521 vdd_d vss_d / DCAP64LVT
XXFILLER_28_606 vdd_d vss_d / DCAP64LVT
XXFILLER_28_670 vdd_d vss_d / DCAP64LVT
XXFILLER_28_734 vdd_d vss_d / DCAP64LVT
XXFILLER_28_798 vdd_d vss_d / DCAP64LVT
XXFILLER_28_920 vdd_d vss_d / DCAP64LVT
XXFILLER_28_984 vdd_d vss_d / DCAP64LVT
XXFILLER_28_1048 vdd_d vss_d / DCAP64LVT
XXFILLER_28_1153 vdd_d vss_d / DCAP64LVT
XXFILLER_28_1249 vdd_d vss_d / DCAP64LVT
XXFILLER_28_1313 vdd_d vss_d / DCAP64LVT
XXFILLER_28_1377 vdd_d vss_d / DCAP64LVT
XXFILLER_28_1441 vdd_d vss_d / DCAP64LVT
XXFILLER_28_1505 vdd_d vss_d / DCAP64LVT
XXFILLER_28_1569 vdd_d vss_d / DCAP64LVT
XXFILLER_28_1633 vdd_d vss_d / DCAP64LVT
XXFILLER_28_1697 vdd_d vss_d / DCAP64LVT
XXFILLER_28_1761 vdd_d vss_d / DCAP64LVT
XXFILLER_28_1825 vdd_d vss_d / DCAP64LVT
XXFILLER_28_1889 vdd_d vss_d / DCAP64LVT
XXFILLER_28_1953 vdd_d vss_d / DCAP64LVT
XXFILLER_28_2017 vdd_d vss_d / DCAP64LVT
XXFILLER_28_2081 vdd_d vss_d / DCAP64LVT
XXFILLER_28_2145 vdd_d vss_d / DCAP64LVT
XXFILLER_28_2209 vdd_d vss_d / DCAP64LVT
XXFILLER_28_2273 vdd_d vss_d / DCAP64LVT
XXFILLER_29_0 vdd_d vss_d / DCAP64LVT
XXFILLER_29_64 vdd_d vss_d / DCAP64LVT
XXFILLER_29_128 vdd_d vss_d / DCAP64LVT
XXFILLER_29_192 vdd_d vss_d / DCAP64LVT
XXFILLER_29_256 vdd_d vss_d / DCAP64LVT
XXFILLER_29_320 vdd_d vss_d / DCAP64LVT
XXFILLER_29_481 vdd_d vss_d / DCAP64LVT
XXFILLER_29_545 vdd_d vss_d / DCAP64LVT
XXFILLER_29_609 vdd_d vss_d / DCAP64LVT
XXFILLER_29_673 vdd_d vss_d / DCAP64LVT
XXFILLER_29_737 vdd_d vss_d / DCAP64LVT
XXFILLER_29_801 vdd_d vss_d / DCAP64LVT
XXFILLER_29_933 vdd_d vss_d / DCAP64LVT
XXFILLER_29_1028 vdd_d vss_d / DCAP64LVT
XXFILLER_29_1092 vdd_d vss_d / DCAP64LVT
XXFILLER_29_1189 vdd_d vss_d / DCAP64LVT
XXFILLER_29_1253 vdd_d vss_d / DCAP64LVT
XXFILLER_29_1343 vdd_d vss_d / DCAP64LVT
XXFILLER_29_1407 vdd_d vss_d / DCAP64LVT
XXFILLER_29_1471 vdd_d vss_d / DCAP64LVT
XXFILLER_29_1535 vdd_d vss_d / DCAP64LVT
XXFILLER_29_1599 vdd_d vss_d / DCAP64LVT
XXFILLER_29_1663 vdd_d vss_d / DCAP64LVT
XXFILLER_29_1727 vdd_d vss_d / DCAP64LVT
XXFILLER_29_1855 vdd_d vss_d / DCAP64LVT
XXFILLER_29_1919 vdd_d vss_d / DCAP64LVT
XXFILLER_29_1983 vdd_d vss_d / DCAP64LVT
XXFILLER_29_2047 vdd_d vss_d / DCAP64LVT
XXFILLER_29_2111 vdd_d vss_d / DCAP64LVT
XXFILLER_29_2175 vdd_d vss_d / DCAP64LVT
XXFILLER_29_2239 vdd_d vss_d / DCAP64LVT
XXFILLER_30_0 vdd_d vss_d / DCAP64LVT
XXFILLER_30_64 vdd_d vss_d / DCAP64LVT
XXFILLER_30_128 vdd_d vss_d / DCAP64LVT
XXFILLER_30_192 vdd_d vss_d / DCAP64LVT
XXFILLER_30_256 vdd_d vss_d / DCAP64LVT
XXFILLER_30_320 vdd_d vss_d / DCAP64LVT
XXFILLER_30_466 vdd_d vss_d / DCAP64LVT
XXFILLER_30_530 vdd_d vss_d / DCAP64LVT
XXFILLER_30_594 vdd_d vss_d / DCAP64LVT
XXFILLER_30_658 vdd_d vss_d / DCAP64LVT
XXFILLER_30_722 vdd_d vss_d / DCAP64LVT
XXFILLER_30_786 vdd_d vss_d / DCAP64LVT
XXFILLER_30_850 vdd_d vss_d / DCAP64LVT
XXFILLER_30_914 vdd_d vss_d / DCAP64LVT
XXFILLER_30_1004 vdd_d vss_d / DCAP64LVT
XXFILLER_30_1068 vdd_d vss_d / DCAP64LVT
XXFILLER_30_1132 vdd_d vss_d / DCAP64LVT
XXFILLER_30_1196 vdd_d vss_d / DCAP64LVT
XXFILLER_30_1260 vdd_d vss_d / DCAP64LVT
XXFILLER_30_1324 vdd_d vss_d / DCAP64LVT
XXFILLER_30_1388 vdd_d vss_d / DCAP64LVT
XXFILLER_30_1452 vdd_d vss_d / DCAP64LVT
XXFILLER_30_1516 vdd_d vss_d / DCAP64LVT
XXFILLER_30_1580 vdd_d vss_d / DCAP64LVT
XXFILLER_30_1644 vdd_d vss_d / DCAP64LVT
XXFILLER_30_1708 vdd_d vss_d / DCAP64LVT
XXFILLER_30_1832 vdd_d vss_d / DCAP64LVT
XXFILLER_30_1896 vdd_d vss_d / DCAP64LVT
XXFILLER_30_1960 vdd_d vss_d / DCAP64LVT
XXFILLER_30_2024 vdd_d vss_d / DCAP64LVT
XXFILLER_30_2088 vdd_d vss_d / DCAP64LVT
XXFILLER_30_2152 vdd_d vss_d / DCAP64LVT
XXFILLER_30_2216 vdd_d vss_d / DCAP64LVT
XXFILLER_30_2280 vdd_d vss_d / DCAP64LVT
XXFILLER_31_0 vdd_d vss_d / DCAP64LVT
XXFILLER_31_64 vdd_d vss_d / DCAP64LVT
XXFILLER_31_128 vdd_d vss_d / DCAP64LVT
XXFILLER_31_192 vdd_d vss_d / DCAP64LVT
XXFILLER_31_256 vdd_d vss_d / DCAP64LVT
XXFILLER_31_320 vdd_d vss_d / DCAP64LVT
XXFILLER_31_518 vdd_d vss_d / DCAP64LVT
XXFILLER_31_582 vdd_d vss_d / DCAP64LVT
XXFILLER_31_646 vdd_d vss_d / DCAP64LVT
XXFILLER_31_710 vdd_d vss_d / DCAP64LVT
XXFILLER_31_818 vdd_d vss_d / DCAP64LVT
XXFILLER_31_882 vdd_d vss_d / DCAP64LVT
XXFILLER_31_946 vdd_d vss_d / DCAP64LVT
XXFILLER_31_1048 vdd_d vss_d / DCAP64LVT
XXFILLER_31_1112 vdd_d vss_d / DCAP64LVT
XXFILLER_31_1176 vdd_d vss_d / DCAP64LVT
XXFILLER_31_1240 vdd_d vss_d / DCAP64LVT
XXFILLER_31_1304 vdd_d vss_d / DCAP64LVT
XXFILLER_31_1368 vdd_d vss_d / DCAP64LVT
XXFILLER_31_1496 vdd_d vss_d / DCAP64LVT
XXFILLER_31_1560 vdd_d vss_d / DCAP64LVT
XXFILLER_31_1624 vdd_d vss_d / DCAP64LVT
XXFILLER_31_1688 vdd_d vss_d / DCAP64LVT
XXFILLER_31_1752 vdd_d vss_d / DCAP64LVT
XXFILLER_31_1892 vdd_d vss_d / DCAP64LVT
XXFILLER_31_1956 vdd_d vss_d / DCAP64LVT
XXFILLER_31_2020 vdd_d vss_d / DCAP64LVT
XXFILLER_31_2084 vdd_d vss_d / DCAP64LVT
XXFILLER_31_2148 vdd_d vss_d / DCAP64LVT
XXFILLER_31_2212 vdd_d vss_d / DCAP64LVT
XXFILLER_31_2276 vdd_d vss_d / DCAP64LVT
XXFILLER_32_0 vdd_d vss_d / DCAP64LVT
XXFILLER_32_64 vdd_d vss_d / DCAP64LVT
XXFILLER_32_128 vdd_d vss_d / DCAP64LVT
XXFILLER_32_192 vdd_d vss_d / DCAP64LVT
XXFILLER_32_256 vdd_d vss_d / DCAP64LVT
XXFILLER_32_320 vdd_d vss_d / DCAP64LVT
XXFILLER_32_428 vdd_d vss_d / DCAP64LVT
XXFILLER_32_492 vdd_d vss_d / DCAP64LVT
XXFILLER_32_556 vdd_d vss_d / DCAP64LVT
XXFILLER_32_620 vdd_d vss_d / DCAP64LVT
XXFILLER_32_684 vdd_d vss_d / DCAP64LVT
XXFILLER_32_806 vdd_d vss_d / DCAP64LVT
XXFILLER_32_870 vdd_d vss_d / DCAP64LVT
XXFILLER_32_998 vdd_d vss_d / DCAP64LVT
XXFILLER_32_1137 vdd_d vss_d / DCAP64LVT
XXFILLER_32_1201 vdd_d vss_d / DCAP64LVT
XXFILLER_32_1265 vdd_d vss_d / DCAP64LVT
XXFILLER_32_1329 vdd_d vss_d / DCAP64LVT
XXFILLER_32_1549 vdd_d vss_d / DCAP64LVT
XXFILLER_32_1613 vdd_d vss_d / DCAP64LVT
XXFILLER_32_1677 vdd_d vss_d / DCAP64LVT
XXFILLER_32_1741 vdd_d vss_d / DCAP64LVT
XXFILLER_32_1862 vdd_d vss_d / DCAP64LVT
XXFILLER_32_1926 vdd_d vss_d / DCAP64LVT
XXFILLER_32_1990 vdd_d vss_d / DCAP64LVT
XXFILLER_32_2054 vdd_d vss_d / DCAP64LVT
XXFILLER_32_2118 vdd_d vss_d / DCAP64LVT
XXFILLER_32_2182 vdd_d vss_d / DCAP64LVT
XXFILLER_32_2246 vdd_d vss_d / DCAP64LVT
XXFILLER_33_0 vdd_d vss_d / DCAP64LVT
XXFILLER_33_64 vdd_d vss_d / DCAP64LVT
XXFILLER_33_128 vdd_d vss_d / DCAP64LVT
XXFILLER_33_192 vdd_d vss_d / DCAP64LVT
XXFILLER_33_256 vdd_d vss_d / DCAP64LVT
XXFILLER_33_320 vdd_d vss_d / DCAP64LVT
XXFILLER_33_478 vdd_d vss_d / DCAP64LVT
XXFILLER_33_542 vdd_d vss_d / DCAP64LVT
XXFILLER_33_606 vdd_d vss_d / DCAP64LVT
XXFILLER_33_670 vdd_d vss_d / DCAP64LVT
XXFILLER_33_734 vdd_d vss_d / DCAP64LVT
XXFILLER_33_798 vdd_d vss_d / DCAP64LVT
XXFILLER_33_862 vdd_d vss_d / DCAP64LVT
XXFILLER_33_967 vdd_d vss_d / DCAP64LVT
XXFILLER_33_1031 vdd_d vss_d / DCAP64LVT
XXFILLER_33_1343 vdd_d vss_d / DCAP64LVT
XXFILLER_33_1495 vdd_d vss_d / DCAP64LVT
XXFILLER_33_1559 vdd_d vss_d / DCAP64LVT
XXFILLER_33_1623 vdd_d vss_d / DCAP64LVT
XXFILLER_33_1687 vdd_d vss_d / DCAP64LVT
XXFILLER_33_1807 vdd_d vss_d / DCAP64LVT
XXFILLER_33_1871 vdd_d vss_d / DCAP64LVT
XXFILLER_33_1935 vdd_d vss_d / DCAP64LVT
XXFILLER_33_1999 vdd_d vss_d / DCAP64LVT
XXFILLER_33_2063 vdd_d vss_d / DCAP64LVT
XXFILLER_33_2127 vdd_d vss_d / DCAP64LVT
XXFILLER_33_2191 vdd_d vss_d / DCAP64LVT
XXFILLER_33_2255 vdd_d vss_d / DCAP64LVT
XXFILLER_34_0 vdd_d vss_d / DCAP64LVT
XXFILLER_34_64 vdd_d vss_d / DCAP64LVT
XXFILLER_34_128 vdd_d vss_d / DCAP64LVT
XXFILLER_34_192 vdd_d vss_d / DCAP64LVT
XXFILLER_34_256 vdd_d vss_d / DCAP64LVT
XXFILLER_34_320 vdd_d vss_d / DCAP64LVT
XXFILLER_34_431 vdd_d vss_d / DCAP64LVT
XXFILLER_34_495 vdd_d vss_d / DCAP64LVT
XXFILLER_34_559 vdd_d vss_d / DCAP64LVT
XXFILLER_34_623 vdd_d vss_d / DCAP64LVT
XXFILLER_34_687 vdd_d vss_d / DCAP64LVT
XXFILLER_34_751 vdd_d vss_d / DCAP64LVT
XXFILLER_34_815 vdd_d vss_d / DCAP64LVT
XXFILLER_34_1241 vdd_d vss_d / DCAP64LVT
XXFILLER_34_1305 vdd_d vss_d / DCAP64LVT
XXFILLER_34_1426 vdd_d vss_d / DCAP64LVT
XXFILLER_34_1567 vdd_d vss_d / DCAP64LVT
XXFILLER_34_1631 vdd_d vss_d / DCAP64LVT
XXFILLER_34_1695 vdd_d vss_d / DCAP64LVT
XXFILLER_34_1759 vdd_d vss_d / DCAP64LVT
XXFILLER_34_1823 vdd_d vss_d / DCAP64LVT
XXFILLER_34_1887 vdd_d vss_d / DCAP64LVT
XXFILLER_34_1951 vdd_d vss_d / DCAP64LVT
XXFILLER_34_2015 vdd_d vss_d / DCAP64LVT
XXFILLER_34_2079 vdd_d vss_d / DCAP64LVT
XXFILLER_34_2143 vdd_d vss_d / DCAP64LVT
XXFILLER_34_2207 vdd_d vss_d / DCAP64LVT
XXFILLER_34_2271 vdd_d vss_d / DCAP64LVT
XXFILLER_35_0 vdd_d vss_d / DCAP64LVT
XXFILLER_35_64 vdd_d vss_d / DCAP64LVT
XXFILLER_35_128 vdd_d vss_d / DCAP64LVT
XXFILLER_35_192 vdd_d vss_d / DCAP64LVT
XXFILLER_35_256 vdd_d vss_d / DCAP64LVT
XXFILLER_35_320 vdd_d vss_d / DCAP64LVT
XXFILLER_35_384 vdd_d vss_d / DCAP64LVT
XXFILLER_35_592 vdd_d vss_d / DCAP64LVT
XXFILLER_35_656 vdd_d vss_d / DCAP64LVT
XXFILLER_35_720 vdd_d vss_d / DCAP64LVT
XXFILLER_35_784 vdd_d vss_d / DCAP64LVT
XXFILLER_35_1096 vdd_d vss_d / DCAP64LVT
XXFILLER_35_1309 vdd_d vss_d / DCAP64LVT
XXFILLER_35_1595 vdd_d vss_d / DCAP64LVT
XXFILLER_35_1659 vdd_d vss_d / DCAP64LVT
XXFILLER_35_1723 vdd_d vss_d / DCAP64LVT
XXFILLER_35_1787 vdd_d vss_d / DCAP64LVT
XXFILLER_35_1851 vdd_d vss_d / DCAP64LVT
XXFILLER_35_1915 vdd_d vss_d / DCAP64LVT
XXFILLER_35_1979 vdd_d vss_d / DCAP64LVT
XXFILLER_35_2043 vdd_d vss_d / DCAP64LVT
XXFILLER_35_2107 vdd_d vss_d / DCAP64LVT
XXFILLER_35_2171 vdd_d vss_d / DCAP64LVT
XXFILLER_35_2235 vdd_d vss_d / DCAP64LVT
XXFILLER_36_0 vdd_d vss_d / DCAP64LVT
XXFILLER_36_64 vdd_d vss_d / DCAP64LVT
XXFILLER_36_128 vdd_d vss_d / DCAP64LVT
XXFILLER_36_192 vdd_d vss_d / DCAP64LVT
XXFILLER_36_256 vdd_d vss_d / DCAP64LVT
XXFILLER_36_320 vdd_d vss_d / DCAP64LVT
XXFILLER_36_419 vdd_d vss_d / DCAP64LVT
XXFILLER_36_483 vdd_d vss_d / DCAP64LVT
XXFILLER_36_547 vdd_d vss_d / DCAP64LVT
XXFILLER_36_611 vdd_d vss_d / DCAP64LVT
XXFILLER_36_675 vdd_d vss_d / DCAP64LVT
XXFILLER_36_1332 vdd_d vss_d / DCAP64LVT
XXFILLER_36_1593 vdd_d vss_d / DCAP64LVT
XXFILLER_36_1657 vdd_d vss_d / DCAP64LVT
XXFILLER_36_1721 vdd_d vss_d / DCAP64LVT
XXFILLER_36_1808 vdd_d vss_d / DCAP64LVT
XXFILLER_36_1892 vdd_d vss_d / DCAP64LVT
XXFILLER_36_1956 vdd_d vss_d / DCAP64LVT
XXFILLER_36_2020 vdd_d vss_d / DCAP64LVT
XXFILLER_36_2084 vdd_d vss_d / DCAP64LVT
XXFILLER_36_2148 vdd_d vss_d / DCAP64LVT
XXFILLER_36_2212 vdd_d vss_d / DCAP64LVT
XXFILLER_36_2276 vdd_d vss_d / DCAP64LVT
XXFILLER_37_0 vdd_d vss_d / DCAP64LVT
XXFILLER_37_64 vdd_d vss_d / DCAP64LVT
XXFILLER_37_128 vdd_d vss_d / DCAP64LVT
XXFILLER_37_192 vdd_d vss_d / DCAP64LVT
XXFILLER_37_256 vdd_d vss_d / DCAP64LVT
XXFILLER_37_320 vdd_d vss_d / DCAP64LVT
XXFILLER_37_546 vdd_d vss_d / DCAP64LVT
XXFILLER_37_610 vdd_d vss_d / DCAP64LVT
XXFILLER_37_674 vdd_d vss_d / DCAP64LVT
XXFILLER_37_973 vdd_d vss_d / DCAP64LVT
XXFILLER_37_1037 vdd_d vss_d / DCAP64LVT
XXFILLER_37_1531 vdd_d vss_d / DCAP64LVT
XXFILLER_37_1692 vdd_d vss_d / DCAP64LVT
XXFILLER_37_1756 vdd_d vss_d / DCAP64LVT
XXFILLER_37_1840 vdd_d vss_d / DCAP64LVT
XXFILLER_37_1931 vdd_d vss_d / DCAP64LVT
XXFILLER_37_1995 vdd_d vss_d / DCAP64LVT
XXFILLER_37_2059 vdd_d vss_d / DCAP64LVT
XXFILLER_37_2123 vdd_d vss_d / DCAP64LVT
XXFILLER_37_2187 vdd_d vss_d / DCAP64LVT
XXFILLER_37_2251 vdd_d vss_d / DCAP64LVT
XXFILLER_38_0 vdd_d vss_d / DCAP64LVT
XXFILLER_38_64 vdd_d vss_d / DCAP64LVT
XXFILLER_38_128 vdd_d vss_d / DCAP64LVT
XXFILLER_38_192 vdd_d vss_d / DCAP64LVT
XXFILLER_38_256 vdd_d vss_d / DCAP64LVT
XXFILLER_38_320 vdd_d vss_d / DCAP64LVT
XXFILLER_38_461 vdd_d vss_d / DCAP64LVT
XXFILLER_38_525 vdd_d vss_d / DCAP64LVT
XXFILLER_38_676 vdd_d vss_d / DCAP64LVT
XXFILLER_38_1125 vdd_d vss_d / DCAP64LVT
XXFILLER_38_1970 vdd_d vss_d / DCAP64LVT
XXFILLER_38_2034 vdd_d vss_d / DCAP64LVT
XXFILLER_38_2098 vdd_d vss_d / DCAP64LVT
XXFILLER_38_2162 vdd_d vss_d / DCAP64LVT
XXFILLER_38_2226 vdd_d vss_d / DCAP64LVT
XXFILLER_39_0 vdd_d vss_d / DCAP64LVT
XXFILLER_39_64 vdd_d vss_d / DCAP64LVT
XXFILLER_39_128 vdd_d vss_d / DCAP64LVT
XXFILLER_39_192 vdd_d vss_d / DCAP64LVT
XXFILLER_39_256 vdd_d vss_d / DCAP64LVT
XXFILLER_39_320 vdd_d vss_d / DCAP64LVT
XXFILLER_39_520 vdd_d vss_d / DCAP64LVT
XXFILLER_39_584 vdd_d vss_d / DCAP64LVT
XXFILLER_39_648 vdd_d vss_d / DCAP64LVT
XXFILLER_39_1656 vdd_d vss_d / DCAP64LVT
XXFILLER_39_1720 vdd_d vss_d / DCAP64LVT
XXFILLER_39_1976 vdd_d vss_d / DCAP64LVT
XXFILLER_39_2040 vdd_d vss_d / DCAP64LVT
XXFILLER_39_2104 vdd_d vss_d / DCAP64LVT
XXFILLER_39_2168 vdd_d vss_d / DCAP64LVT
XXFILLER_39_2232 vdd_d vss_d / DCAP64LVT
XXFILLER_40_0 vdd_d vss_d / DCAP64LVT
XXFILLER_40_64 vdd_d vss_d / DCAP64LVT
XXFILLER_40_128 vdd_d vss_d / DCAP64LVT
XXFILLER_40_192 vdd_d vss_d / DCAP64LVT
XXFILLER_40_256 vdd_d vss_d / DCAP64LVT
XXFILLER_40_320 vdd_d vss_d / DCAP64LVT
XXFILLER_40_625 vdd_d vss_d / DCAP64LVT
XXFILLER_40_815 vdd_d vss_d / DCAP64LVT
XXFILLER_40_1691 vdd_d vss_d / DCAP64LVT
XXFILLER_40_1997 vdd_d vss_d / DCAP64LVT
XXFILLER_40_2061 vdd_d vss_d / DCAP64LVT
XXFILLER_40_2125 vdd_d vss_d / DCAP64LVT
XXFILLER_40_2189 vdd_d vss_d / DCAP64LVT
XXFILLER_40_2253 vdd_d vss_d / DCAP64LVT
XXFILLER_41_0 vdd_d vss_d / DCAP64LVT
XXFILLER_41_64 vdd_d vss_d / DCAP64LVT
XXFILLER_41_128 vdd_d vss_d / DCAP64LVT
XXFILLER_41_192 vdd_d vss_d / DCAP64LVT
XXFILLER_41_256 vdd_d vss_d / DCAP64LVT
XXFILLER_41_320 vdd_d vss_d / DCAP64LVT
XXFILLER_41_512 vdd_d vss_d / DCAP64LVT
XXFILLER_41_576 vdd_d vss_d / DCAP64LVT
XXFILLER_41_640 vdd_d vss_d / DCAP64LVT
XXFILLER_41_704 vdd_d vss_d / DCAP64LVT
XXFILLER_41_1622 vdd_d vss_d / DCAP64LVT
XXFILLER_41_1739 vdd_d vss_d / DCAP64LVT
XXFILLER_41_1987 vdd_d vss_d / DCAP64LVT
XXFILLER_41_2051 vdd_d vss_d / DCAP64LVT
XXFILLER_41_2115 vdd_d vss_d / DCAP64LVT
XXFILLER_41_2179 vdd_d vss_d / DCAP64LVT
XXFILLER_41_2243 vdd_d vss_d / DCAP64LVT
XXFILLER_42_0 vdd_d vss_d / DCAP64LVT
XXFILLER_42_64 vdd_d vss_d / DCAP64LVT
XXFILLER_42_128 vdd_d vss_d / DCAP64LVT
XXFILLER_42_192 vdd_d vss_d / DCAP64LVT
XXFILLER_42_256 vdd_d vss_d / DCAP64LVT
XXFILLER_42_320 vdd_d vss_d / DCAP64LVT
XXFILLER_42_486 vdd_d vss_d / DCAP64LVT
XXFILLER_42_604 vdd_d vss_d / DCAP64LVT
XXFILLER_42_1017 vdd_d vss_d / DCAP64LVT
XXFILLER_42_1701 vdd_d vss_d / DCAP64LVT
XXFILLER_42_1819 vdd_d vss_d / DCAP64LVT
XXFILLER_42_2040 vdd_d vss_d / DCAP64LVT
XXFILLER_42_2104 vdd_d vss_d / DCAP64LVT
XXFILLER_42_2168 vdd_d vss_d / DCAP64LVT
XXFILLER_42_2232 vdd_d vss_d / DCAP64LVT
XXFILLER_43_0 vdd_d vss_d / DCAP64LVT
XXFILLER_43_64 vdd_d vss_d / DCAP64LVT
XXFILLER_43_128 vdd_d vss_d / DCAP64LVT
XXFILLER_43_192 vdd_d vss_d / DCAP64LVT
XXFILLER_43_256 vdd_d vss_d / DCAP64LVT
XXFILLER_43_320 vdd_d vss_d / DCAP64LVT
XXFILLER_43_429 vdd_d vss_d / DCAP64LVT
XXFILLER_43_515 vdd_d vss_d / DCAP64LVT
XXFILLER_43_579 vdd_d vss_d / DCAP64LVT
XXFILLER_43_643 vdd_d vss_d / DCAP64LVT
XXFILLER_43_956 vdd_d vss_d / DCAP64LVT
XXFILLER_43_1020 vdd_d vss_d / DCAP64LVT
XXFILLER_43_1681 vdd_d vss_d / DCAP64LVT
XXFILLER_43_1986 vdd_d vss_d / DCAP64LVT
XXFILLER_43_2050 vdd_d vss_d / DCAP64LVT
XXFILLER_43_2114 vdd_d vss_d / DCAP64LVT
XXFILLER_43_2178 vdd_d vss_d / DCAP64LVT
XXFILLER_43_2242 vdd_d vss_d / DCAP64LVT
XXFILLER_44_0 vdd_d vss_d / DCAP64LVT
XXFILLER_44_64 vdd_d vss_d / DCAP64LVT
XXFILLER_44_128 vdd_d vss_d / DCAP64LVT
XXFILLER_44_192 vdd_d vss_d / DCAP64LVT
XXFILLER_44_256 vdd_d vss_d / DCAP64LVT
XXFILLER_44_494 vdd_d vss_d / DCAP64LVT
XXFILLER_44_558 vdd_d vss_d / DCAP64LVT
XXFILLER_44_622 vdd_d vss_d / DCAP64LVT
XXFILLER_44_1753 vdd_d vss_d / DCAP64LVT
XXFILLER_44_1946 vdd_d vss_d / DCAP64LVT
XXFILLER_44_2010 vdd_d vss_d / DCAP64LVT
XXFILLER_44_2074 vdd_d vss_d / DCAP64LVT
XXFILLER_44_2138 vdd_d vss_d / DCAP64LVT
XXFILLER_44_2202 vdd_d vss_d / DCAP64LVT
XXFILLER_44_2266 vdd_d vss_d / DCAP64LVT
XXFILLER_45_0 vdd_d vss_d / DCAP64LVT
XXFILLER_45_64 vdd_d vss_d / DCAP64LVT
XXFILLER_45_128 vdd_d vss_d / DCAP64LVT
XXFILLER_45_192 vdd_d vss_d / DCAP64LVT
XXFILLER_45_256 vdd_d vss_d / DCAP64LVT
XXFILLER_45_320 vdd_d vss_d / DCAP64LVT
XXFILLER_45_384 vdd_d vss_d / DCAP64LVT
XXFILLER_45_448 vdd_d vss_d / DCAP64LVT
XXFILLER_45_512 vdd_d vss_d / DCAP64LVT
XXFILLER_45_576 vdd_d vss_d / DCAP64LVT
XXFILLER_45_640 vdd_d vss_d / DCAP64LVT
XXFILLER_45_736 vdd_d vss_d / DCAP64LVT
XXFILLER_45_860 vdd_d vss_d / DCAP64LVT
XXFILLER_45_938 vdd_d vss_d / DCAP64LVT
XXFILLER_45_1016 vdd_d vss_d / DCAP64LVT
XXFILLER_45_1080 vdd_d vss_d / DCAP64LVT
XXFILLER_45_1144 vdd_d vss_d / DCAP64LVT
XXFILLER_45_1208 vdd_d vss_d / DCAP64LVT
XXFILLER_45_1272 vdd_d vss_d / DCAP64LVT
XXFILLER_45_1336 vdd_d vss_d / DCAP64LVT
XXFILLER_45_1400 vdd_d vss_d / DCAP64LVT
XXFILLER_45_1464 vdd_d vss_d / DCAP64LVT
XXFILLER_45_1654 vdd_d vss_d / DCAP64LVT
XXFILLER_45_1718 vdd_d vss_d / DCAP64LVT
XXFILLER_45_1782 vdd_d vss_d / DCAP64LVT
XXFILLER_45_1907 vdd_d vss_d / DCAP64LVT
XXFILLER_45_1971 vdd_d vss_d / DCAP64LVT
XXFILLER_45_2035 vdd_d vss_d / DCAP64LVT
XXFILLER_45_2099 vdd_d vss_d / DCAP64LVT
XXFILLER_45_2163 vdd_d vss_d / DCAP64LVT
XXFILLER_45_2227 vdd_d vss_d / DCAP64LVT
XXFILLER_46_0 vdd_d vss_d / DCAP64LVT
XXFILLER_46_64 vdd_d vss_d / DCAP64LVT
XXFILLER_46_128 vdd_d vss_d / DCAP64LVT
XXFILLER_46_192 vdd_d vss_d / DCAP64LVT
XXFILLER_46_256 vdd_d vss_d / DCAP64LVT
XXFILLER_46_320 vdd_d vss_d / DCAP64LVT
XXFILLER_46_384 vdd_d vss_d / DCAP64LVT
XXFILLER_46_448 vdd_d vss_d / DCAP64LVT
XXFILLER_46_512 vdd_d vss_d / DCAP64LVT
XXFILLER_46_576 vdd_d vss_d / DCAP64LVT
XXFILLER_46_640 vdd_d vss_d / DCAP64LVT
XXFILLER_46_704 vdd_d vss_d / DCAP64LVT
XXFILLER_46_768 vdd_d vss_d / DCAP64LVT
XXFILLER_46_832 vdd_d vss_d / DCAP64LVT
XXFILLER_46_910 vdd_d vss_d / DCAP64LVT
XXFILLER_46_974 vdd_d vss_d / DCAP64LVT
XXFILLER_46_1038 vdd_d vss_d / DCAP64LVT
XXFILLER_46_1102 vdd_d vss_d / DCAP64LVT
XXFILLER_46_1166 vdd_d vss_d / DCAP64LVT
XXFILLER_46_1230 vdd_d vss_d / DCAP64LVT
XXFILLER_46_1294 vdd_d vss_d / DCAP64LVT
XXFILLER_46_1410 vdd_d vss_d / DCAP64LVT
XXFILLER_46_1474 vdd_d vss_d / DCAP64LVT
XXFILLER_46_1552 vdd_d vss_d / DCAP64LVT
XXFILLER_46_1616 vdd_d vss_d / DCAP64LVT
XXFILLER_46_1713 vdd_d vss_d / DCAP64LVT
XXFILLER_46_1777 vdd_d vss_d / DCAP64LVT
XXFILLER_46_1841 vdd_d vss_d / DCAP64LVT
XXFILLER_46_1983 vdd_d vss_d / DCAP64LVT
XXFILLER_46_2047 vdd_d vss_d / DCAP64LVT
XXFILLER_46_2111 vdd_d vss_d / DCAP64LVT
XXFILLER_46_2175 vdd_d vss_d / DCAP64LVT
XXFILLER_46_2239 vdd_d vss_d / DCAP64LVT
XXFILLER_47_0 vdd_d vss_d / DCAP64LVT
XXFILLER_47_64 vdd_d vss_d / DCAP64LVT
XXFILLER_47_128 vdd_d vss_d / DCAP64LVT
XXFILLER_47_192 vdd_d vss_d / DCAP64LVT
XXFILLER_47_256 vdd_d vss_d / DCAP64LVT
XXFILLER_47_320 vdd_d vss_d / DCAP64LVT
XXFILLER_47_384 vdd_d vss_d / DCAP64LVT
XXFILLER_47_448 vdd_d vss_d / DCAP64LVT
XXFILLER_47_512 vdd_d vss_d / DCAP64LVT
XXFILLER_47_576 vdd_d vss_d / DCAP64LVT
XXFILLER_47_680 vdd_d vss_d / DCAP64LVT
XXFILLER_47_744 vdd_d vss_d / DCAP64LVT
XXFILLER_47_808 vdd_d vss_d / DCAP64LVT
XXFILLER_47_872 vdd_d vss_d / DCAP64LVT
XXFILLER_47_936 vdd_d vss_d / DCAP64LVT
XXFILLER_47_1000 vdd_d vss_d / DCAP64LVT
XXFILLER_47_1064 vdd_d vss_d / DCAP64LVT
XXFILLER_47_1128 vdd_d vss_d / DCAP64LVT
XXFILLER_47_1192 vdd_d vss_d / DCAP64LVT
XXFILLER_47_1256 vdd_d vss_d / DCAP64LVT
XXFILLER_47_1320 vdd_d vss_d / DCAP64LVT
XXFILLER_47_1384 vdd_d vss_d / DCAP64LVT
XXFILLER_47_1448 vdd_d vss_d / DCAP64LVT
XXFILLER_47_1512 vdd_d vss_d / DCAP64LVT
XXFILLER_47_1576 vdd_d vss_d / DCAP64LVT
XXFILLER_47_1640 vdd_d vss_d / DCAP64LVT
XXFILLER_47_1704 vdd_d vss_d / DCAP64LVT
XXFILLER_47_1768 vdd_d vss_d / DCAP64LVT
XXFILLER_47_1832 vdd_d vss_d / DCAP64LVT
XXFILLER_47_1896 vdd_d vss_d / DCAP64LVT
XXFILLER_47_1960 vdd_d vss_d / DCAP64LVT
XXFILLER_47_2024 vdd_d vss_d / DCAP64LVT
XXFILLER_47_2088 vdd_d vss_d / DCAP64LVT
XXFILLER_47_2152 vdd_d vss_d / DCAP64LVT
XXFILLER_47_2216 vdd_d vss_d / DCAP64LVT
XXFILLER_47_2280 vdd_d vss_d / DCAP64LVT
XXFILLER_48_0 vdd_d vss_d / DCAP64LVT
XXFILLER_48_103 vdd_d vss_d / DCAP64LVT
XXFILLER_48_167 vdd_d vss_d / DCAP64LVT
XXFILLER_48_231 vdd_d vss_d / DCAP64LVT
XXFILLER_48_295 vdd_d vss_d / DCAP64LVT
XXFILLER_48_370 vdd_d vss_d / DCAP64LVT
XXFILLER_48_434 vdd_d vss_d / DCAP64LVT
XXFILLER_48_498 vdd_d vss_d / DCAP64LVT
XXFILLER_48_562 vdd_d vss_d / DCAP64LVT
XXFILLER_48_626 vdd_d vss_d / DCAP64LVT
XXFILLER_48_690 vdd_d vss_d / DCAP64LVT
XXFILLER_48_754 vdd_d vss_d / DCAP64LVT
XXFILLER_48_818 vdd_d vss_d / DCAP64LVT
XXFILLER_48_925 vdd_d vss_d / DCAP64LVT
XXFILLER_48_989 vdd_d vss_d / DCAP64LVT
XXFILLER_48_1053 vdd_d vss_d / DCAP64LVT
XXFILLER_48_1117 vdd_d vss_d / DCAP64LVT
XXFILLER_48_1181 vdd_d vss_d / DCAP64LVT
XXFILLER_48_1245 vdd_d vss_d / DCAP64LVT
XXFILLER_48_1309 vdd_d vss_d / DCAP64LVT
XXFILLER_48_1373 vdd_d vss_d / DCAP64LVT
XXFILLER_48_1437 vdd_d vss_d / DCAP64LVT
XXFILLER_48_1501 vdd_d vss_d / DCAP64LVT
XXFILLER_48_1565 vdd_d vss_d / DCAP64LVT
XXFILLER_48_1629 vdd_d vss_d / DCAP64LVT
XXFILLER_48_1693 vdd_d vss_d / DCAP64LVT
XXFILLER_48_1757 vdd_d vss_d / DCAP64LVT
XXFILLER_48_1821 vdd_d vss_d / DCAP64LVT
XXFILLER_48_1885 vdd_d vss_d / DCAP64LVT
XXFILLER_48_1949 vdd_d vss_d / DCAP64LVT
XXFILLER_48_2013 vdd_d vss_d / DCAP64LVT
XXFILLER_48_2077 vdd_d vss_d / DCAP64LVT
XXFILLER_48_2141 vdd_d vss_d / DCAP64LVT
XXFILLER_48_2271 vdd_d vss_d / DCAP64LVT
XXFILLER_49_0 vdd_d vss_d / DCAP64LVT
XXFILLER_49_64 vdd_d vss_d / DCAP64LVT
XXFILLER_49_128 vdd_d vss_d / DCAP64LVT
XXFILLER_49_192 vdd_d vss_d / DCAP64LVT
XXFILLER_49_256 vdd_d vss_d / DCAP64LVT
XXFILLER_49_320 vdd_d vss_d / DCAP64LVT
XXFILLER_49_423 vdd_d vss_d / DCAP64LVT
XXFILLER_49_487 vdd_d vss_d / DCAP64LVT
XXFILLER_49_551 vdd_d vss_d / DCAP64LVT
XXFILLER_49_615 vdd_d vss_d / DCAP64LVT
XXFILLER_49_679 vdd_d vss_d / DCAP64LVT
XXFILLER_49_743 vdd_d vss_d / DCAP64LVT
XXFILLER_49_807 vdd_d vss_d / DCAP64LVT
XXFILLER_49_871 vdd_d vss_d / DCAP64LVT
XXFILLER_49_935 vdd_d vss_d / DCAP64LVT
XXFILLER_49_999 vdd_d vss_d / DCAP64LVT
XXFILLER_49_1063 vdd_d vss_d / DCAP64LVT
XXFILLER_49_1127 vdd_d vss_d / DCAP64LVT
XXFILLER_49_1191 vdd_d vss_d / DCAP64LVT
XXFILLER_49_1255 vdd_d vss_d / DCAP64LVT
XXFILLER_49_1319 vdd_d vss_d / DCAP64LVT
XXFILLER_49_1383 vdd_d vss_d / DCAP64LVT
XXFILLER_49_1521 vdd_d vss_d / DCAP64LVT
XXFILLER_49_1585 vdd_d vss_d / DCAP64LVT
XXFILLER_49_1649 vdd_d vss_d / DCAP64LVT
XXFILLER_49_1713 vdd_d vss_d / DCAP64LVT
XXFILLER_49_1777 vdd_d vss_d / DCAP64LVT
XXFILLER_49_1841 vdd_d vss_d / DCAP64LVT
XXFILLER_49_1905 vdd_d vss_d / DCAP64LVT
XXFILLER_49_1969 vdd_d vss_d / DCAP64LVT
XXFILLER_49_2033 vdd_d vss_d / DCAP64LVT
XXFILLER_49_2097 vdd_d vss_d / DCAP64LVT
XXFILLER_49_2161 vdd_d vss_d / DCAP64LVT
XXFILLER_49_2225 vdd_d vss_d / DCAP64LVT
XXFILLER_50_0 vdd_d vss_d / DCAP64LVT
XXFILLER_50_64 vdd_d vss_d / DCAP64LVT
XXFILLER_50_128 vdd_d vss_d / DCAP64LVT
XXFILLER_50_192 vdd_d vss_d / DCAP64LVT
XXFILLER_50_256 vdd_d vss_d / DCAP64LVT
XXFILLER_50_320 vdd_d vss_d / DCAP64LVT
XXFILLER_50_443 vdd_d vss_d / DCAP64LVT
XXFILLER_50_507 vdd_d vss_d / DCAP64LVT
XXFILLER_50_571 vdd_d vss_d / DCAP64LVT
XXFILLER_50_635 vdd_d vss_d / DCAP64LVT
XXFILLER_50_699 vdd_d vss_d / DCAP64LVT
XXFILLER_50_829 vdd_d vss_d / DCAP64LVT
XXFILLER_50_893 vdd_d vss_d / DCAP64LVT
XXFILLER_50_957 vdd_d vss_d / DCAP64LVT
XXFILLER_50_1021 vdd_d vss_d / DCAP64LVT
XXFILLER_50_1085 vdd_d vss_d / DCAP64LVT
XXFILLER_50_1149 vdd_d vss_d / DCAP64LVT
XXFILLER_50_1213 vdd_d vss_d / DCAP64LVT
XXFILLER_50_1277 vdd_d vss_d / DCAP64LVT
XXFILLER_50_1341 vdd_d vss_d / DCAP64LVT
XXFILLER_50_1405 vdd_d vss_d / DCAP64LVT
XXFILLER_50_1521 vdd_d vss_d / DCAP64LVT
XXFILLER_50_1585 vdd_d vss_d / DCAP64LVT
XXFILLER_50_1649 vdd_d vss_d / DCAP64LVT
XXFILLER_50_1770 vdd_d vss_d / DCAP64LVT
XXFILLER_50_1834 vdd_d vss_d / DCAP64LVT
XXFILLER_50_1950 vdd_d vss_d / DCAP64LVT
XXFILLER_50_2014 vdd_d vss_d / DCAP64LVT
XXFILLER_50_2078 vdd_d vss_d / DCAP64LVT
XXFILLER_50_2142 vdd_d vss_d / DCAP64LVT
XXFILLER_50_2206 vdd_d vss_d / DCAP64LVT
XXFILLER_50_2270 vdd_d vss_d / DCAP64LVT
XXFILLER_51_0 vdd_d vss_d / DCAP64LVT
XXFILLER_51_64 vdd_d vss_d / DCAP64LVT
XXFILLER_51_128 vdd_d vss_d / DCAP64LVT
XXFILLER_51_192 vdd_d vss_d / DCAP64LVT
XXFILLER_51_256 vdd_d vss_d / DCAP64LVT
XXFILLER_51_320 vdd_d vss_d / DCAP64LVT
XXFILLER_51_384 vdd_d vss_d / DCAP64LVT
XXFILLER_51_448 vdd_d vss_d / DCAP64LVT
XXFILLER_51_512 vdd_d vss_d / DCAP64LVT
XXFILLER_51_576 vdd_d vss_d / DCAP64LVT
XXFILLER_51_640 vdd_d vss_d / DCAP64LVT
XXFILLER_51_704 vdd_d vss_d / DCAP64LVT
XXFILLER_51_768 vdd_d vss_d / DCAP64LVT
XXFILLER_51_832 vdd_d vss_d / DCAP64LVT
XXFILLER_51_896 vdd_d vss_d / DCAP64LVT
XXFILLER_51_960 vdd_d vss_d / DCAP64LVT
XXFILLER_51_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_51_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_51_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_51_1293 vdd_d vss_d / DCAP64LVT
XXFILLER_51_1357 vdd_d vss_d / DCAP64LVT
XXFILLER_51_1421 vdd_d vss_d / DCAP64LVT
XXFILLER_51_1485 vdd_d vss_d / DCAP64LVT
XXFILLER_51_1549 vdd_d vss_d / DCAP64LVT
XXFILLER_51_1613 vdd_d vss_d / DCAP64LVT
XXFILLER_51_1677 vdd_d vss_d / DCAP64LVT
XXFILLER_51_1741 vdd_d vss_d / DCAP64LVT
XXFILLER_51_1805 vdd_d vss_d / DCAP64LVT
XXFILLER_51_1869 vdd_d vss_d / DCAP64LVT
XXFILLER_51_1933 vdd_d vss_d / DCAP64LVT
XXFILLER_51_1997 vdd_d vss_d / DCAP64LVT
XXFILLER_51_2061 vdd_d vss_d / DCAP64LVT
XXFILLER_51_2125 vdd_d vss_d / DCAP64LVT
XXFILLER_51_2189 vdd_d vss_d / DCAP64LVT
XXFILLER_51_2253 vdd_d vss_d / DCAP64LVT
XXFILLER_52_0 vdd_d vss_d / DCAP64LVT
XXFILLER_52_64 vdd_d vss_d / DCAP64LVT
XXFILLER_52_128 vdd_d vss_d / DCAP64LVT
XXFILLER_52_192 vdd_d vss_d / DCAP64LVT
XXFILLER_52_256 vdd_d vss_d / DCAP64LVT
XXFILLER_52_320 vdd_d vss_d / DCAP64LVT
XXFILLER_52_384 vdd_d vss_d / DCAP64LVT
XXFILLER_52_448 vdd_d vss_d / DCAP64LVT
XXFILLER_52_512 vdd_d vss_d / DCAP64LVT
XXFILLER_52_576 vdd_d vss_d / DCAP64LVT
XXFILLER_52_640 vdd_d vss_d / DCAP64LVT
XXFILLER_52_704 vdd_d vss_d / DCAP64LVT
XXFILLER_52_768 vdd_d vss_d / DCAP64LVT
XXFILLER_52_832 vdd_d vss_d / DCAP64LVT
XXFILLER_52_896 vdd_d vss_d / DCAP64LVT
XXFILLER_52_960 vdd_d vss_d / DCAP64LVT
XXFILLER_52_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_52_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_52_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_52_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_52_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_52_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_52_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_52_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_52_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_52_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_52_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_52_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_52_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_52_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_52_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_52_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_52_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_52_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_52_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_52_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_53_0 vdd_d vss_d / DCAP64LVT
XXFILLER_53_64 vdd_d vss_d / DCAP64LVT
XXFILLER_53_128 vdd_d vss_d / DCAP64LVT
XXFILLER_53_192 vdd_d vss_d / DCAP64LVT
XXFILLER_53_256 vdd_d vss_d / DCAP64LVT
XXFILLER_53_320 vdd_d vss_d / DCAP64LVT
XXFILLER_53_384 vdd_d vss_d / DCAP64LVT
XXFILLER_53_448 vdd_d vss_d / DCAP64LVT
XXFILLER_53_512 vdd_d vss_d / DCAP64LVT
XXFILLER_53_576 vdd_d vss_d / DCAP64LVT
XXFILLER_53_640 vdd_d vss_d / DCAP64LVT
XXFILLER_53_704 vdd_d vss_d / DCAP64LVT
XXFILLER_53_768 vdd_d vss_d / DCAP64LVT
XXFILLER_53_832 vdd_d vss_d / DCAP64LVT
XXFILLER_53_896 vdd_d vss_d / DCAP64LVT
XXFILLER_53_960 vdd_d vss_d / DCAP64LVT
XXFILLER_53_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_53_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_53_1232 vdd_d vss_d / DCAP64LVT
XXFILLER_53_1296 vdd_d vss_d / DCAP64LVT
XXFILLER_53_1360 vdd_d vss_d / DCAP64LVT
XXFILLER_53_1424 vdd_d vss_d / DCAP64LVT
XXFILLER_53_1488 vdd_d vss_d / DCAP64LVT
XXFILLER_53_1552 vdd_d vss_d / DCAP64LVT
XXFILLER_53_1616 vdd_d vss_d / DCAP64LVT
XXFILLER_53_1680 vdd_d vss_d / DCAP64LVT
XXFILLER_53_1744 vdd_d vss_d / DCAP64LVT
XXFILLER_53_1808 vdd_d vss_d / DCAP64LVT
XXFILLER_53_1872 vdd_d vss_d / DCAP64LVT
XXFILLER_53_1936 vdd_d vss_d / DCAP64LVT
XXFILLER_53_2000 vdd_d vss_d / DCAP64LVT
XXFILLER_53_2064 vdd_d vss_d / DCAP64LVT
XXFILLER_53_2128 vdd_d vss_d / DCAP64LVT
XXFILLER_53_2192 vdd_d vss_d / DCAP64LVT
XXFILLER_53_2256 vdd_d vss_d / DCAP64LVT
XXFILLER_54_0 vdd_d vss_d / DCAP64LVT
XXFILLER_54_64 vdd_d vss_d / DCAP64LVT
XXFILLER_54_128 vdd_d vss_d / DCAP64LVT
XXFILLER_54_192 vdd_d vss_d / DCAP64LVT
XXFILLER_54_256 vdd_d vss_d / DCAP64LVT
XXFILLER_54_320 vdd_d vss_d / DCAP64LVT
XXFILLER_54_384 vdd_d vss_d / DCAP64LVT
XXFILLER_54_448 vdd_d vss_d / DCAP64LVT
XXFILLER_54_512 vdd_d vss_d / DCAP64LVT
XXFILLER_54_576 vdd_d vss_d / DCAP64LVT
XXFILLER_54_640 vdd_d vss_d / DCAP64LVT
XXFILLER_54_704 vdd_d vss_d / DCAP64LVT
XXFILLER_54_935 vdd_d vss_d / DCAP64LVT
XXFILLER_54_999 vdd_d vss_d / DCAP64LVT
XXFILLER_54_1063 vdd_d vss_d / DCAP64LVT
XXFILLER_54_1127 vdd_d vss_d / DCAP64LVT
XXFILLER_54_1191 vdd_d vss_d / DCAP64LVT
XXFILLER_54_1255 vdd_d vss_d / DCAP64LVT
XXFILLER_54_1319 vdd_d vss_d / DCAP64LVT
XXFILLER_54_1383 vdd_d vss_d / DCAP64LVT
XXFILLER_54_1447 vdd_d vss_d / DCAP64LVT
XXFILLER_54_1511 vdd_d vss_d / DCAP64LVT
XXFILLER_54_1575 vdd_d vss_d / DCAP64LVT
XXFILLER_54_1639 vdd_d vss_d / DCAP64LVT
XXFILLER_54_1703 vdd_d vss_d / DCAP64LVT
XXFILLER_54_1767 vdd_d vss_d / DCAP64LVT
XXFILLER_54_1831 vdd_d vss_d / DCAP64LVT
XXFILLER_54_1965 vdd_d vss_d / DCAP64LVT
XXFILLER_54_2029 vdd_d vss_d / DCAP64LVT
XXFILLER_54_2093 vdd_d vss_d / DCAP64LVT
XXFILLER_54_2157 vdd_d vss_d / DCAP64LVT
XXFILLER_54_2221 vdd_d vss_d / DCAP64LVT
XXFILLER_54_2285 vdd_d vss_d / DCAP64LVT
XXFILLER_55_0 vdd_d vss_d / DCAP64LVT
XXFILLER_55_64 vdd_d vss_d / DCAP64LVT
XXFILLER_55_128 vdd_d vss_d / DCAP64LVT
XXFILLER_55_192 vdd_d vss_d / DCAP64LVT
XXFILLER_55_256 vdd_d vss_d / DCAP64LVT
XXFILLER_55_320 vdd_d vss_d / DCAP64LVT
XXFILLER_55_437 vdd_d vss_d / DCAP64LVT
XXFILLER_55_501 vdd_d vss_d / DCAP64LVT
XXFILLER_55_565 vdd_d vss_d / DCAP64LVT
XXFILLER_55_629 vdd_d vss_d / DCAP64LVT
XXFILLER_55_693 vdd_d vss_d / DCAP64LVT
XXFILLER_55_757 vdd_d vss_d / DCAP64LVT
XXFILLER_55_821 vdd_d vss_d / DCAP64LVT
XXFILLER_55_944 vdd_d vss_d / DCAP64LVT
XXFILLER_55_1008 vdd_d vss_d / DCAP64LVT
XXFILLER_55_1072 vdd_d vss_d / DCAP64LVT
XXFILLER_55_1136 vdd_d vss_d / DCAP64LVT
XXFILLER_55_1200 vdd_d vss_d / DCAP64LVT
XXFILLER_55_1264 vdd_d vss_d / DCAP64LVT
XXFILLER_55_1328 vdd_d vss_d / DCAP64LVT
XXFILLER_55_1392 vdd_d vss_d / DCAP64LVT
XXFILLER_55_1456 vdd_d vss_d / DCAP64LVT
XXFILLER_55_1520 vdd_d vss_d / DCAP64LVT
XXFILLER_55_1584 vdd_d vss_d / DCAP64LVT
XXFILLER_55_1648 vdd_d vss_d / DCAP64LVT
XXFILLER_55_1712 vdd_d vss_d / DCAP64LVT
XXFILLER_55_1776 vdd_d vss_d / DCAP64LVT
XXFILLER_55_1840 vdd_d vss_d / DCAP64LVT
XXFILLER_55_1978 vdd_d vss_d / DCAP64LVT
XXFILLER_55_2042 vdd_d vss_d / DCAP64LVT
XXFILLER_55_2106 vdd_d vss_d / DCAP64LVT
XXFILLER_55_2170 vdd_d vss_d / DCAP64LVT
XXFILLER_55_2234 vdd_d vss_d / DCAP64LVT
XXFILLER_56_0 vdd_d vss_d / DCAP64LVT
XXFILLER_56_64 vdd_d vss_d / DCAP64LVT
XXFILLER_56_128 vdd_d vss_d / DCAP64LVT
XXFILLER_56_192 vdd_d vss_d / DCAP64LVT
XXFILLER_56_587 vdd_d vss_d / DCAP64LVT
XXFILLER_56_651 vdd_d vss_d / DCAP64LVT
XXFILLER_56_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_56_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_56_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_56_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_56_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_56_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_56_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_56_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_57_0 vdd_d vss_d / DCAP64LVT
XXFILLER_57_64 vdd_d vss_d / DCAP64LVT
XXFILLER_57_128 vdd_d vss_d / DCAP64LVT
XXFILLER_57_192 vdd_d vss_d / DCAP64LVT
XXFILLER_57_587 vdd_d vss_d / DCAP64LVT
XXFILLER_57_651 vdd_d vss_d / DCAP64LVT
XXFILLER_57_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_57_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_57_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_57_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_57_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_57_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_57_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_58_0 vdd_d vss_d / DCAP64LVT
XXFILLER_58_64 vdd_d vss_d / DCAP64LVT
XXFILLER_58_128 vdd_d vss_d / DCAP64LVT
XXFILLER_58_192 vdd_d vss_d / DCAP64LVT
XXFILLER_58_587 vdd_d vss_d / DCAP64LVT
XXFILLER_58_651 vdd_d vss_d / DCAP64LVT
XXFILLER_58_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_58_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_58_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_58_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_58_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_58_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_58_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_58_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_59_0 vdd_d vss_d / DCAP64LVT
XXFILLER_59_64 vdd_d vss_d / DCAP64LVT
XXFILLER_59_128 vdd_d vss_d / DCAP64LVT
XXFILLER_59_192 vdd_d vss_d / DCAP64LVT
XXFILLER_59_587 vdd_d vss_d / DCAP64LVT
XXFILLER_59_651 vdd_d vss_d / DCAP64LVT
XXFILLER_59_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_59_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_59_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_59_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_59_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_59_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_59_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_59_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_60_0 vdd_d vss_d / DCAP64LVT
XXFILLER_60_64 vdd_d vss_d / DCAP64LVT
XXFILLER_60_128 vdd_d vss_d / DCAP64LVT
XXFILLER_60_192 vdd_d vss_d / DCAP64LVT
XXFILLER_60_587 vdd_d vss_d / DCAP64LVT
XXFILLER_60_651 vdd_d vss_d / DCAP64LVT
XXFILLER_60_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_60_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_60_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_60_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_60_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_60_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_60_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_60_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_61_0 vdd_d vss_d / DCAP64LVT
XXFILLER_61_64 vdd_d vss_d / DCAP64LVT
XXFILLER_61_128 vdd_d vss_d / DCAP64LVT
XXFILLER_61_192 vdd_d vss_d / DCAP64LVT
XXFILLER_61_587 vdd_d vss_d / DCAP64LVT
XXFILLER_61_651 vdd_d vss_d / DCAP64LVT
XXFILLER_61_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_61_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_61_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_61_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_61_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_61_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_61_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_61_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_62_0 vdd_d vss_d / DCAP64LVT
XXFILLER_62_64 vdd_d vss_d / DCAP64LVT
XXFILLER_62_128 vdd_d vss_d / DCAP64LVT
XXFILLER_62_192 vdd_d vss_d / DCAP64LVT
XXFILLER_62_587 vdd_d vss_d / DCAP64LVT
XXFILLER_62_651 vdd_d vss_d / DCAP64LVT
XXFILLER_62_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_62_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_62_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_62_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_62_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_62_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_62_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_62_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_63_0 vdd_d vss_d / DCAP64LVT
XXFILLER_63_64 vdd_d vss_d / DCAP64LVT
XXFILLER_63_128 vdd_d vss_d / DCAP64LVT
XXFILLER_63_192 vdd_d vss_d / DCAP64LVT
XXFILLER_63_587 vdd_d vss_d / DCAP64LVT
XXFILLER_63_651 vdd_d vss_d / DCAP64LVT
XXFILLER_63_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_63_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_63_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_63_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_63_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_63_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_63_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_63_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_64_0 vdd_d vss_d / DCAP64LVT
XXFILLER_64_64 vdd_d vss_d / DCAP64LVT
XXFILLER_64_128 vdd_d vss_d / DCAP64LVT
XXFILLER_64_192 vdd_d vss_d / DCAP64LVT
XXFILLER_64_587 vdd_d vss_d / DCAP64LVT
XXFILLER_64_651 vdd_d vss_d / DCAP64LVT
XXFILLER_64_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_64_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_64_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_64_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_64_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_64_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_64_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_64_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_65_0 vdd_d vss_d / DCAP64LVT
XXFILLER_65_64 vdd_d vss_d / DCAP64LVT
XXFILLER_65_128 vdd_d vss_d / DCAP64LVT
XXFILLER_65_192 vdd_d vss_d / DCAP64LVT
XXFILLER_65_587 vdd_d vss_d / DCAP64LVT
XXFILLER_65_651 vdd_d vss_d / DCAP64LVT
XXFILLER_65_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_65_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_65_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_65_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_65_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_65_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_65_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_65_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_66_0 vdd_d vss_d / DCAP64LVT
XXFILLER_66_64 vdd_d vss_d / DCAP64LVT
XXFILLER_66_128 vdd_d vss_d / DCAP64LVT
XXFILLER_66_192 vdd_d vss_d / DCAP64LVT
XXFILLER_66_587 vdd_d vss_d / DCAP64LVT
XXFILLER_66_651 vdd_d vss_d / DCAP64LVT
XXFILLER_66_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_66_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_66_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_66_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_66_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_66_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_66_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_66_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_67_0 vdd_d vss_d / DCAP64LVT
XXFILLER_67_64 vdd_d vss_d / DCAP64LVT
XXFILLER_67_128 vdd_d vss_d / DCAP64LVT
XXFILLER_67_192 vdd_d vss_d / DCAP64LVT
XXFILLER_67_587 vdd_d vss_d / DCAP64LVT
XXFILLER_67_651 vdd_d vss_d / DCAP64LVT
XXFILLER_67_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_67_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_67_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_67_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_67_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_67_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_67_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_67_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_68_0 vdd_d vss_d / DCAP64LVT
XXFILLER_68_64 vdd_d vss_d / DCAP64LVT
XXFILLER_68_128 vdd_d vss_d / DCAP64LVT
XXFILLER_68_192 vdd_d vss_d / DCAP64LVT
XXFILLER_68_587 vdd_d vss_d / DCAP64LVT
XXFILLER_68_651 vdd_d vss_d / DCAP64LVT
XXFILLER_68_1093 vdd_d vss_d / DCAP64LVT
XXFILLER_68_1157 vdd_d vss_d / DCAP64LVT
XXFILLER_68_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_68_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_68_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_68_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_68_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_68_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_69_0 vdd_d vss_d / DCAP64LVT
XXFILLER_69_64 vdd_d vss_d / DCAP64LVT
XXFILLER_69_128 vdd_d vss_d / DCAP64LVT
XXFILLER_69_587 vdd_d vss_d / DCAP64LVT
XXFILLER_69_651 vdd_d vss_d / DCAP64LVT
XXFILLER_69_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_69_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_69_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_69_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_69_2103 vdd_d vss_d / DCAP64LVT
XXFILLER_69_2167 vdd_d vss_d / DCAP64LVT
XXFILLER_69_2231 vdd_d vss_d / DCAP64LVT
XXFILLER_70_0 vdd_d vss_d / DCAP64LVT
XXFILLER_70_64 vdd_d vss_d / DCAP64LVT
XXFILLER_70_128 vdd_d vss_d / DCAP64LVT
XXFILLER_70_192 vdd_d vss_d / DCAP64LVT
XXFILLER_70_587 vdd_d vss_d / DCAP64LVT
XXFILLER_70_651 vdd_d vss_d / DCAP64LVT
XXFILLER_70_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_70_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_70_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_70_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_70_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_70_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_70_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_70_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_71_0 vdd_d vss_d / DCAP64LVT
XXFILLER_71_64 vdd_d vss_d / DCAP64LVT
XXFILLER_71_128 vdd_d vss_d / DCAP64LVT
XXFILLER_71_192 vdd_d vss_d / DCAP64LVT
XXFILLER_71_587 vdd_d vss_d / DCAP64LVT
XXFILLER_71_651 vdd_d vss_d / DCAP64LVT
XXFILLER_71_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_71_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_71_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_71_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_71_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_71_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_71_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_71_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_72_0 vdd_d vss_d / DCAP64LVT
XXFILLER_72_64 vdd_d vss_d / DCAP64LVT
XXFILLER_72_128 vdd_d vss_d / DCAP64LVT
XXFILLER_72_192 vdd_d vss_d / DCAP64LVT
XXFILLER_72_587 vdd_d vss_d / DCAP64LVT
XXFILLER_72_651 vdd_d vss_d / DCAP64LVT
XXFILLER_72_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_72_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_72_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_72_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_72_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_72_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_72_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_73_0 vdd_d vss_d / DCAP64LVT
XXFILLER_73_64 vdd_d vss_d / DCAP64LVT
XXFILLER_73_128 vdd_d vss_d / DCAP64LVT
XXFILLER_73_587 vdd_d vss_d / DCAP64LVT
XXFILLER_73_651 vdd_d vss_d / DCAP64LVT
XXFILLER_73_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_73_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_73_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_73_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_73_2122 vdd_d vss_d / DCAP64LVT
XXFILLER_73_2186 vdd_d vss_d / DCAP64LVT
XXFILLER_73_2250 vdd_d vss_d / DCAP64LVT
XXFILLER_74_0 vdd_d vss_d / DCAP64LVT
XXFILLER_74_64 vdd_d vss_d / DCAP64LVT
XXFILLER_74_128 vdd_d vss_d / DCAP64LVT
XXFILLER_74_192 vdd_d vss_d / DCAP64LVT
XXFILLER_74_587 vdd_d vss_d / DCAP64LVT
XXFILLER_74_651 vdd_d vss_d / DCAP64LVT
XXFILLER_74_1137 vdd_d vss_d / DCAP64LVT
XXFILLER_74_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_74_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_74_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_74_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_74_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_74_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_75_0 vdd_d vss_d / DCAP64LVT
XXFILLER_75_64 vdd_d vss_d / DCAP64LVT
XXFILLER_75_128 vdd_d vss_d / DCAP64LVT
XXFILLER_75_192 vdd_d vss_d / DCAP64LVT
XXFILLER_75_587 vdd_d vss_d / DCAP64LVT
XXFILLER_75_651 vdd_d vss_d / DCAP64LVT
XXFILLER_75_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_75_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_75_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_75_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_75_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_75_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_75_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_75_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_76_0 vdd_d vss_d / DCAP64LVT
XXFILLER_76_64 vdd_d vss_d / DCAP64LVT
XXFILLER_76_128 vdd_d vss_d / DCAP64LVT
XXFILLER_76_587 vdd_d vss_d / DCAP64LVT
XXFILLER_76_651 vdd_d vss_d / DCAP64LVT
XXFILLER_76_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_76_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_76_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_76_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_76_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_76_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_76_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_76_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_77_0 vdd_d vss_d / DCAP64LVT
XXFILLER_77_64 vdd_d vss_d / DCAP64LVT
XXFILLER_77_128 vdd_d vss_d / DCAP64LVT
XXFILLER_77_192 vdd_d vss_d / DCAP64LVT
XXFILLER_77_587 vdd_d vss_d / DCAP64LVT
XXFILLER_77_651 vdd_d vss_d / DCAP64LVT
XXFILLER_77_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_77_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_77_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_77_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_77_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_77_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_77_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_78_0 vdd_d vss_d / DCAP64LVT
XXFILLER_78_64 vdd_d vss_d / DCAP64LVT
XXFILLER_78_128 vdd_d vss_d / DCAP64LVT
XXFILLER_78_192 vdd_d vss_d / DCAP64LVT
XXFILLER_78_587 vdd_d vss_d / DCAP64LVT
XXFILLER_78_651 vdd_d vss_d / DCAP64LVT
XXFILLER_78_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_78_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_78_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_78_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_78_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_78_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_78_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_78_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_79_0 vdd_d vss_d / DCAP64LVT
XXFILLER_79_64 vdd_d vss_d / DCAP64LVT
XXFILLER_79_128 vdd_d vss_d / DCAP64LVT
XXFILLER_79_192 vdd_d vss_d / DCAP64LVT
XXFILLER_79_587 vdd_d vss_d / DCAP64LVT
XXFILLER_79_651 vdd_d vss_d / DCAP64LVT
XXFILLER_79_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_79_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_79_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_79_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_79_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_79_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_79_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_79_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_80_0 vdd_d vss_d / DCAP64LVT
XXFILLER_80_64 vdd_d vss_d / DCAP64LVT
XXFILLER_80_128 vdd_d vss_d / DCAP64LVT
XXFILLER_80_192 vdd_d vss_d / DCAP64LVT
XXFILLER_80_587 vdd_d vss_d / DCAP64LVT
XXFILLER_80_651 vdd_d vss_d / DCAP64LVT
XXFILLER_80_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_80_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_80_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_80_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_80_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_80_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_80_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_80_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_81_0 vdd_d vss_d / DCAP64LVT
XXFILLER_81_64 vdd_d vss_d / DCAP64LVT
XXFILLER_81_128 vdd_d vss_d / DCAP64LVT
XXFILLER_81_192 vdd_d vss_d / DCAP64LVT
XXFILLER_81_587 vdd_d vss_d / DCAP64LVT
XXFILLER_81_651 vdd_d vss_d / DCAP64LVT
XXFILLER_81_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_81_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_81_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_81_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_81_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_81_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_81_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_81_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_82_0 vdd_d vss_d / DCAP64LVT
XXFILLER_82_64 vdd_d vss_d / DCAP64LVT
XXFILLER_82_128 vdd_d vss_d / DCAP64LVT
XXFILLER_82_192 vdd_d vss_d / DCAP64LVT
XXFILLER_82_587 vdd_d vss_d / DCAP64LVT
XXFILLER_82_651 vdd_d vss_d / DCAP64LVT
XXFILLER_82_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_82_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_82_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_82_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_82_2096 vdd_d vss_d / DCAP64LVT
XXFILLER_82_2160 vdd_d vss_d / DCAP64LVT
XXFILLER_82_2224 vdd_d vss_d / DCAP64LVT
XXFILLER_83_0 vdd_d vss_d / DCAP64LVT
XXFILLER_83_64 vdd_d vss_d / DCAP64LVT
XXFILLER_83_128 vdd_d vss_d / DCAP64LVT
XXFILLER_83_587 vdd_d vss_d / DCAP64LVT
XXFILLER_83_651 vdd_d vss_d / DCAP64LVT
XXFILLER_83_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_83_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_83_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_83_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_83_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_83_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_83_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_83_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_84_0 vdd_d vss_d / DCAP64LVT
XXFILLER_84_64 vdd_d vss_d / DCAP64LVT
XXFILLER_84_128 vdd_d vss_d / DCAP64LVT
XXFILLER_84_192 vdd_d vss_d / DCAP64LVT
XXFILLER_84_587 vdd_d vss_d / DCAP64LVT
XXFILLER_84_651 vdd_d vss_d / DCAP64LVT
XXFILLER_84_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_84_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_84_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_84_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_84_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_84_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_84_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_84_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_85_0 vdd_d vss_d / DCAP64LVT
XXFILLER_85_64 vdd_d vss_d / DCAP64LVT
XXFILLER_85_128 vdd_d vss_d / DCAP64LVT
XXFILLER_85_192 vdd_d vss_d / DCAP64LVT
XXFILLER_85_587 vdd_d vss_d / DCAP64LVT
XXFILLER_85_651 vdd_d vss_d / DCAP64LVT
XXFILLER_85_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_85_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_85_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_85_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_85_2096 vdd_d vss_d / DCAP64LVT
XXFILLER_85_2160 vdd_d vss_d / DCAP64LVT
XXFILLER_85_2224 vdd_d vss_d / DCAP64LVT
XXFILLER_86_0 vdd_d vss_d / DCAP64LVT
XXFILLER_86_64 vdd_d vss_d / DCAP64LVT
XXFILLER_86_128 vdd_d vss_d / DCAP64LVT
XXFILLER_86_192 vdd_d vss_d / DCAP64LVT
XXFILLER_86_587 vdd_d vss_d / DCAP64LVT
XXFILLER_86_651 vdd_d vss_d / DCAP64LVT
XXFILLER_86_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_86_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_86_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_86_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_86_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_86_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_86_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_86_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_87_0 vdd_d vss_d / DCAP64LVT
XXFILLER_87_64 vdd_d vss_d / DCAP64LVT
XXFILLER_87_128 vdd_d vss_d / DCAP64LVT
XXFILLER_87_192 vdd_d vss_d / DCAP64LVT
XXFILLER_87_587 vdd_d vss_d / DCAP64LVT
XXFILLER_87_651 vdd_d vss_d / DCAP64LVT
XXFILLER_87_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_87_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_87_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_87_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_87_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_87_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_87_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_87_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_88_0 vdd_d vss_d / DCAP64LVT
XXFILLER_88_64 vdd_d vss_d / DCAP64LVT
XXFILLER_88_128 vdd_d vss_d / DCAP64LVT
XXFILLER_88_192 vdd_d vss_d / DCAP64LVT
XXFILLER_88_587 vdd_d vss_d / DCAP64LVT
XXFILLER_88_651 vdd_d vss_d / DCAP64LVT
XXFILLER_88_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_88_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_88_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_88_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_88_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_88_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_88_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_88_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_89_0 vdd_d vss_d / DCAP64LVT
XXFILLER_89_64 vdd_d vss_d / DCAP64LVT
XXFILLER_89_128 vdd_d vss_d / DCAP64LVT
XXFILLER_89_192 vdd_d vss_d / DCAP64LVT
XXFILLER_89_587 vdd_d vss_d / DCAP64LVT
XXFILLER_89_651 vdd_d vss_d / DCAP64LVT
XXFILLER_89_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_89_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_89_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_89_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_89_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_89_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_89_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_89_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_90_0 vdd_d vss_d / DCAP64LVT
XXFILLER_90_64 vdd_d vss_d / DCAP64LVT
XXFILLER_90_128 vdd_d vss_d / DCAP64LVT
XXFILLER_90_192 vdd_d vss_d / DCAP64LVT
XXFILLER_90_587 vdd_d vss_d / DCAP64LVT
XXFILLER_90_651 vdd_d vss_d / DCAP64LVT
XXFILLER_90_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_90_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_90_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_90_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_90_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_90_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_90_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_90_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_91_0 vdd_d vss_d / DCAP64LVT
XXFILLER_91_64 vdd_d vss_d / DCAP64LVT
XXFILLER_91_128 vdd_d vss_d / DCAP64LVT
XXFILLER_91_192 vdd_d vss_d / DCAP64LVT
XXFILLER_91_587 vdd_d vss_d / DCAP64LVT
XXFILLER_91_651 vdd_d vss_d / DCAP64LVT
XXFILLER_91_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_91_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_91_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_91_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_91_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_91_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_91_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_91_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_92_0 vdd_d vss_d / DCAP64LVT
XXFILLER_92_64 vdd_d vss_d / DCAP64LVT
XXFILLER_92_128 vdd_d vss_d / DCAP64LVT
XXFILLER_92_192 vdd_d vss_d / DCAP64LVT
XXFILLER_92_587 vdd_d vss_d / DCAP64LVT
XXFILLER_92_651 vdd_d vss_d / DCAP64LVT
XXFILLER_92_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_92_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_92_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_92_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_92_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_92_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_92_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_92_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_93_0 vdd_d vss_d / DCAP64LVT
XXFILLER_93_64 vdd_d vss_d / DCAP64LVT
XXFILLER_93_128 vdd_d vss_d / DCAP64LVT
XXFILLER_93_192 vdd_d vss_d / DCAP64LVT
XXFILLER_93_587 vdd_d vss_d / DCAP64LVT
XXFILLER_93_651 vdd_d vss_d / DCAP64LVT
XXFILLER_93_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_93_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_93_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_93_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_93_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_93_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_93_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_93_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_94_0 vdd_d vss_d / DCAP64LVT
XXFILLER_94_64 vdd_d vss_d / DCAP64LVT
XXFILLER_94_128 vdd_d vss_d / DCAP64LVT
XXFILLER_94_192 vdd_d vss_d / DCAP64LVT
XXFILLER_94_635 vdd_d vss_d / DCAP64LVT
XXFILLER_94_699 vdd_d vss_d / DCAP64LVT
XXFILLER_94_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_94_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_94_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_94_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_94_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_94_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_94_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_94_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_95_0 vdd_d vss_d / DCAP64LVT
XXFILLER_95_64 vdd_d vss_d / DCAP64LVT
XXFILLER_95_128 vdd_d vss_d / DCAP64LVT
XXFILLER_95_192 vdd_d vss_d / DCAP64LVT
XXFILLER_95_256 vdd_d vss_d / DCAP64LVT
XXFILLER_95_320 vdd_d vss_d / DCAP64LVT
XXFILLER_95_475 vdd_d vss_d / DCAP64LVT
XXFILLER_95_539 vdd_d vss_d / DCAP64LVT
XXFILLER_95_603 vdd_d vss_d / DCAP64LVT
XXFILLER_95_667 vdd_d vss_d / DCAP64LVT
XXFILLER_95_731 vdd_d vss_d / DCAP64LVT
XXFILLER_95_795 vdd_d vss_d / DCAP64LVT
XXFILLER_95_859 vdd_d vss_d / DCAP64LVT
XXFILLER_95_988 vdd_d vss_d / DCAP64LVT
XXFILLER_95_1052 vdd_d vss_d / DCAP64LVT
XXFILLER_95_1116 vdd_d vss_d / DCAP64LVT
XXFILLER_95_1180 vdd_d vss_d / DCAP64LVT
XXFILLER_95_1244 vdd_d vss_d / DCAP64LVT
XXFILLER_95_1308 vdd_d vss_d / DCAP64LVT
XXFILLER_95_1451 vdd_d vss_d / DCAP64LVT
XXFILLER_95_1515 vdd_d vss_d / DCAP64LVT
XXFILLER_95_1579 vdd_d vss_d / DCAP64LVT
XXFILLER_95_1643 vdd_d vss_d / DCAP64LVT
XXFILLER_95_1707 vdd_d vss_d / DCAP64LVT
XXFILLER_95_1771 vdd_d vss_d / DCAP64LVT
XXFILLER_95_1899 vdd_d vss_d / DCAP64LVT
XXFILLER_95_1963 vdd_d vss_d / DCAP64LVT
XXFILLER_95_2027 vdd_d vss_d / DCAP64LVT
XXFILLER_95_2091 vdd_d vss_d / DCAP64LVT
XXFILLER_95_2155 vdd_d vss_d / DCAP64LVT
XXFILLER_95_2219 vdd_d vss_d / DCAP64LVT
XXFILLER_95_2283 vdd_d vss_d / DCAP64LVT
XXFILLER_96_0 vdd_d vss_d / DCAP64LVT
XXFILLER_96_64 vdd_d vss_d / DCAP64LVT
XXFILLER_96_128 vdd_d vss_d / DCAP64LVT
XXFILLER_96_192 vdd_d vss_d / DCAP64LVT
XXFILLER_96_256 vdd_d vss_d / DCAP64LVT
XXFILLER_96_459 vdd_d vss_d / DCAP64LVT
XXFILLER_96_523 vdd_d vss_d / DCAP64LVT
XXFILLER_96_587 vdd_d vss_d / DCAP64LVT
XXFILLER_96_651 vdd_d vss_d / DCAP64LVT
XXFILLER_96_715 vdd_d vss_d / DCAP64LVT
XXFILLER_96_779 vdd_d vss_d / DCAP64LVT
XXFILLER_96_843 vdd_d vss_d / DCAP64LVT
XXFILLER_96_907 vdd_d vss_d / DCAP64LVT
XXFILLER_96_971 vdd_d vss_d / DCAP64LVT
XXFILLER_96_1035 vdd_d vss_d / DCAP64LVT
XXFILLER_96_1099 vdd_d vss_d / DCAP64LVT
XXFILLER_96_1163 vdd_d vss_d / DCAP64LVT
XXFILLER_96_1227 vdd_d vss_d / DCAP64LVT
XXFILLER_96_1291 vdd_d vss_d / DCAP64LVT
XXFILLER_96_1460 vdd_d vss_d / DCAP64LVT
XXFILLER_96_1524 vdd_d vss_d / DCAP64LVT
XXFILLER_96_1588 vdd_d vss_d / DCAP64LVT
XXFILLER_96_1652 vdd_d vss_d / DCAP64LVT
XXFILLER_96_1716 vdd_d vss_d / DCAP64LVT
XXFILLER_96_1780 vdd_d vss_d / DCAP64LVT
XXFILLER_96_1844 vdd_d vss_d / DCAP64LVT
XXFILLER_96_1908 vdd_d vss_d / DCAP64LVT
XXFILLER_96_1972 vdd_d vss_d / DCAP64LVT
XXFILLER_96_2036 vdd_d vss_d / DCAP64LVT
XXFILLER_96_2100 vdd_d vss_d / DCAP64LVT
XXFILLER_96_2164 vdd_d vss_d / DCAP64LVT
XXFILLER_96_2228 vdd_d vss_d / DCAP64LVT
XXFILLER_97_0 vdd_d vss_d / DCAP64LVT
XXFILLER_97_64 vdd_d vss_d / DCAP64LVT
XXFILLER_97_128 vdd_d vss_d / DCAP64LVT
XXFILLER_97_192 vdd_d vss_d / DCAP64LVT
XXFILLER_97_256 vdd_d vss_d / DCAP64LVT
XXFILLER_97_385 vdd_d vss_d / DCAP64LVT
XXFILLER_97_470 vdd_d vss_d / DCAP64LVT
XXFILLER_97_534 vdd_d vss_d / DCAP64LVT
XXFILLER_97_598 vdd_d vss_d / DCAP64LVT
XXFILLER_97_662 vdd_d vss_d / DCAP64LVT
XXFILLER_97_726 vdd_d vss_d / DCAP64LVT
XXFILLER_97_790 vdd_d vss_d / DCAP64LVT
XXFILLER_97_854 vdd_d vss_d / DCAP64LVT
XXFILLER_97_918 vdd_d vss_d / DCAP64LVT
XXFILLER_97_982 vdd_d vss_d / DCAP64LVT
XXFILLER_97_1046 vdd_d vss_d / DCAP64LVT
XXFILLER_97_1110 vdd_d vss_d / DCAP64LVT
XXFILLER_97_1174 vdd_d vss_d / DCAP64LVT
XXFILLER_97_1238 vdd_d vss_d / DCAP64LVT
XXFILLER_97_1302 vdd_d vss_d / DCAP64LVT
XXFILLER_97_1366 vdd_d vss_d / DCAP64LVT
XXFILLER_97_1462 vdd_d vss_d / DCAP64LVT
XXFILLER_97_1526 vdd_d vss_d / DCAP64LVT
XXFILLER_97_1590 vdd_d vss_d / DCAP64LVT
XXFILLER_97_1654 vdd_d vss_d / DCAP64LVT
XXFILLER_97_1718 vdd_d vss_d / DCAP64LVT
XXFILLER_97_1782 vdd_d vss_d / DCAP64LVT
XXFILLER_97_1846 vdd_d vss_d / DCAP64LVT
XXFILLER_97_1910 vdd_d vss_d / DCAP64LVT
XXFILLER_97_1974 vdd_d vss_d / DCAP64LVT
XXFILLER_97_2038 vdd_d vss_d / DCAP64LVT
XXFILLER_97_2102 vdd_d vss_d / DCAP64LVT
XXFILLER_97_2166 vdd_d vss_d / DCAP64LVT
XXFILLER_97_2230 vdd_d vss_d / DCAP64LVT
XXFILLER_98_0 vdd_d vss_d / DCAP64LVT
XXFILLER_98_64 vdd_d vss_d / DCAP64LVT
XXFILLER_98_128 vdd_d vss_d / DCAP64LVT
XXFILLER_98_192 vdd_d vss_d / DCAP64LVT
XXFILLER_98_256 vdd_d vss_d / DCAP64LVT
XXFILLER_98_320 vdd_d vss_d / DCAP64LVT
XXFILLER_98_421 vdd_d vss_d / DCAP64LVT
XXFILLER_98_485 vdd_d vss_d / DCAP64LVT
XXFILLER_98_549 vdd_d vss_d / DCAP64LVT
XXFILLER_98_613 vdd_d vss_d / DCAP64LVT
XXFILLER_98_677 vdd_d vss_d / DCAP64LVT
XXFILLER_98_741 vdd_d vss_d / DCAP64LVT
XXFILLER_98_805 vdd_d vss_d / DCAP64LVT
XXFILLER_98_869 vdd_d vss_d / DCAP64LVT
XXFILLER_98_933 vdd_d vss_d / DCAP64LVT
XXFILLER_98_997 vdd_d vss_d / DCAP64LVT
XXFILLER_98_1061 vdd_d vss_d / DCAP64LVT
XXFILLER_98_1125 vdd_d vss_d / DCAP64LVT
XXFILLER_98_1189 vdd_d vss_d / DCAP64LVT
XXFILLER_98_1253 vdd_d vss_d / DCAP64LVT
XXFILLER_98_1317 vdd_d vss_d / DCAP64LVT
XXFILLER_98_1381 vdd_d vss_d / DCAP64LVT
XXFILLER_98_1445 vdd_d vss_d / DCAP64LVT
XXFILLER_98_1545 vdd_d vss_d / DCAP64LVT
XXFILLER_98_1628 vdd_d vss_d / DCAP64LVT
XXFILLER_98_1692 vdd_d vss_d / DCAP64LVT
XXFILLER_98_1812 vdd_d vss_d / DCAP64LVT
XXFILLER_98_1876 vdd_d vss_d / DCAP64LVT
XXFILLER_98_1940 vdd_d vss_d / DCAP64LVT
XXFILLER_98_2004 vdd_d vss_d / DCAP64LVT
XXFILLER_98_2068 vdd_d vss_d / DCAP64LVT
XXFILLER_98_2132 vdd_d vss_d / DCAP64LVT
XXFILLER_98_2196 vdd_d vss_d / DCAP64LVT
XXFILLER_98_2260 vdd_d vss_d / DCAP64LVT
XXFILLER_99_0 vdd_d vss_d / DCAP64LVT
XXFILLER_99_64 vdd_d vss_d / DCAP64LVT
XXFILLER_99_128 vdd_d vss_d / DCAP64LVT
XXFILLER_99_192 vdd_d vss_d / DCAP64LVT
XXFILLER_99_256 vdd_d vss_d / DCAP64LVT
XXFILLER_99_320 vdd_d vss_d / DCAP64LVT
XXFILLER_99_384 vdd_d vss_d / DCAP64LVT
XXFILLER_99_448 vdd_d vss_d / DCAP64LVT
XXFILLER_99_512 vdd_d vss_d / DCAP64LVT
XXFILLER_99_576 vdd_d vss_d / DCAP64LVT
XXFILLER_99_640 vdd_d vss_d / DCAP64LVT
XXFILLER_99_704 vdd_d vss_d / DCAP64LVT
XXFILLER_99_768 vdd_d vss_d / DCAP64LVT
XXFILLER_99_832 vdd_d vss_d / DCAP64LVT
XXFILLER_99_896 vdd_d vss_d / DCAP64LVT
XXFILLER_99_990 vdd_d vss_d / DCAP64LVT
XXFILLER_99_1054 vdd_d vss_d / DCAP64LVT
XXFILLER_99_1118 vdd_d vss_d / DCAP64LVT
XXFILLER_99_1182 vdd_d vss_d / DCAP64LVT
XXFILLER_99_1246 vdd_d vss_d / DCAP64LVT
XXFILLER_99_1310 vdd_d vss_d / DCAP64LVT
XXFILLER_99_1426 vdd_d vss_d / DCAP64LVT
XXFILLER_99_1490 vdd_d vss_d / DCAP64LVT
XXFILLER_99_1554 vdd_d vss_d / DCAP64LVT
XXFILLER_99_1618 vdd_d vss_d / DCAP64LVT
XXFILLER_99_1682 vdd_d vss_d / DCAP64LVT
XXFILLER_99_1746 vdd_d vss_d / DCAP64LVT
XXFILLER_99_1810 vdd_d vss_d / DCAP64LVT
XXFILLER_99_1928 vdd_d vss_d / DCAP64LVT
XXFILLER_99_1992 vdd_d vss_d / DCAP64LVT
XXFILLER_99_2056 vdd_d vss_d / DCAP64LVT
XXFILLER_99_2120 vdd_d vss_d / DCAP64LVT
XXFILLER_99_2184 vdd_d vss_d / DCAP64LVT
XXFILLER_99_2248 vdd_d vss_d / DCAP64LVT
XXFILLER_100_0 vdd_d vss_d / DCAP64LVT
XXFILLER_100_64 vdd_d vss_d / DCAP64LVT
XXFILLER_100_128 vdd_d vss_d / DCAP64LVT
XXFILLER_100_192 vdd_d vss_d / DCAP64LVT
XXFILLER_100_256 vdd_d vss_d / DCAP64LVT
XXFILLER_100_320 vdd_d vss_d / DCAP64LVT
XXFILLER_100_384 vdd_d vss_d / DCAP64LVT
XXFILLER_100_448 vdd_d vss_d / DCAP64LVT
XXFILLER_100_512 vdd_d vss_d / DCAP64LVT
XXFILLER_100_576 vdd_d vss_d / DCAP64LVT
XXFILLER_100_640 vdd_d vss_d / DCAP64LVT
XXFILLER_100_704 vdd_d vss_d / DCAP64LVT
XXFILLER_100_768 vdd_d vss_d / DCAP64LVT
XXFILLER_100_832 vdd_d vss_d / DCAP64LVT
XXFILLER_100_896 vdd_d vss_d / DCAP64LVT
XXFILLER_100_960 vdd_d vss_d / DCAP64LVT
XXFILLER_100_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_100_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_100_1208 vdd_d vss_d / DCAP64LVT
XXFILLER_100_1272 vdd_d vss_d / DCAP64LVT
XXFILLER_100_1336 vdd_d vss_d / DCAP64LVT
XXFILLER_100_1400 vdd_d vss_d / DCAP64LVT
XXFILLER_100_1464 vdd_d vss_d / DCAP64LVT
XXFILLER_100_1528 vdd_d vss_d / DCAP64LVT
XXFILLER_100_1592 vdd_d vss_d / DCAP64LVT
XXFILLER_100_1656 vdd_d vss_d / DCAP64LVT
XXFILLER_100_1720 vdd_d vss_d / DCAP64LVT
XXFILLER_100_1784 vdd_d vss_d / DCAP64LVT
XXFILLER_100_1848 vdd_d vss_d / DCAP64LVT
XXFILLER_100_1912 vdd_d vss_d / DCAP64LVT
XXFILLER_100_1976 vdd_d vss_d / DCAP64LVT
XXFILLER_100_2040 vdd_d vss_d / DCAP64LVT
XXFILLER_100_2104 vdd_d vss_d / DCAP64LVT
XXFILLER_100_2168 vdd_d vss_d / DCAP64LVT
XXFILLER_100_2232 vdd_d vss_d / DCAP64LVT
XXFILLER_101_0 vdd_d vss_d / DCAP64LVT
XXFILLER_101_64 vdd_d vss_d / DCAP64LVT
XXFILLER_101_128 vdd_d vss_d / DCAP64LVT
XXFILLER_101_192 vdd_d vss_d / DCAP64LVT
XXFILLER_101_256 vdd_d vss_d / DCAP64LVT
XXFILLER_101_320 vdd_d vss_d / DCAP64LVT
XXFILLER_101_384 vdd_d vss_d / DCAP64LVT
XXFILLER_101_448 vdd_d vss_d / DCAP64LVT
XXFILLER_101_512 vdd_d vss_d / DCAP64LVT
XXFILLER_101_576 vdd_d vss_d / DCAP64LVT
XXFILLER_101_640 vdd_d vss_d / DCAP64LVT
XXFILLER_101_704 vdd_d vss_d / DCAP64LVT
XXFILLER_101_768 vdd_d vss_d / DCAP64LVT
XXFILLER_101_832 vdd_d vss_d / DCAP64LVT
XXFILLER_101_896 vdd_d vss_d / DCAP64LVT
XXFILLER_101_960 vdd_d vss_d / DCAP64LVT
XXFILLER_101_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_101_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_101_1213 vdd_d vss_d / DCAP64LVT
XXFILLER_101_1277 vdd_d vss_d / DCAP64LVT
XXFILLER_101_1341 vdd_d vss_d / DCAP64LVT
XXFILLER_101_1405 vdd_d vss_d / DCAP64LVT
XXFILLER_101_1469 vdd_d vss_d / DCAP64LVT
XXFILLER_101_1533 vdd_d vss_d / DCAP64LVT
XXFILLER_101_1597 vdd_d vss_d / DCAP64LVT
XXFILLER_101_1661 vdd_d vss_d / DCAP64LVT
XXFILLER_101_1725 vdd_d vss_d / DCAP64LVT
XXFILLER_101_1789 vdd_d vss_d / DCAP64LVT
XXFILLER_101_1853 vdd_d vss_d / DCAP64LVT
XXFILLER_101_2036 vdd_d vss_d / DCAP64LVT
XXFILLER_101_2100 vdd_d vss_d / DCAP64LVT
XXFILLER_101_2164 vdd_d vss_d / DCAP64LVT
XXFILLER_101_2228 vdd_d vss_d / DCAP64LVT
XXFILLER_102_0 vdd_d vss_d / DCAP64LVT
XXFILLER_102_64 vdd_d vss_d / DCAP64LVT
XXFILLER_102_128 vdd_d vss_d / DCAP64LVT
XXFILLER_102_192 vdd_d vss_d / DCAP64LVT
XXFILLER_102_256 vdd_d vss_d / DCAP64LVT
XXFILLER_102_320 vdd_d vss_d / DCAP64LVT
XXFILLER_102_384 vdd_d vss_d / DCAP64LVT
XXFILLER_102_448 vdd_d vss_d / DCAP64LVT
XXFILLER_102_512 vdd_d vss_d / DCAP64LVT
XXFILLER_102_576 vdd_d vss_d / DCAP64LVT
XXFILLER_102_688 vdd_d vss_d / DCAP64LVT
XXFILLER_102_752 vdd_d vss_d / DCAP64LVT
XXFILLER_102_816 vdd_d vss_d / DCAP64LVT
XXFILLER_102_880 vdd_d vss_d / DCAP64LVT
XXFILLER_102_944 vdd_d vss_d / DCAP64LVT
XXFILLER_102_1070 vdd_d vss_d / DCAP64LVT
XXFILLER_102_1198 vdd_d vss_d / DCAP64LVT
XXFILLER_102_1348 vdd_d vss_d / DCAP64LVT
XXFILLER_102_1412 vdd_d vss_d / DCAP64LVT
XXFILLER_102_1476 vdd_d vss_d / DCAP64LVT
XXFILLER_102_1540 vdd_d vss_d / DCAP64LVT
XXFILLER_102_1604 vdd_d vss_d / DCAP64LVT
XXFILLER_102_1668 vdd_d vss_d / DCAP64LVT
XXFILLER_102_1732 vdd_d vss_d / DCAP64LVT
XXFILLER_102_1796 vdd_d vss_d / DCAP64LVT
XXFILLER_102_1860 vdd_d vss_d / DCAP64LVT
XXFILLER_102_1924 vdd_d vss_d / DCAP64LVT
XXFILLER_102_1988 vdd_d vss_d / DCAP64LVT
XXFILLER_102_2052 vdd_d vss_d / DCAP64LVT
XXFILLER_102_2116 vdd_d vss_d / DCAP64LVT
XXFILLER_102_2180 vdd_d vss_d / DCAP64LVT
XXFILLER_102_2244 vdd_d vss_d / DCAP64LVT
XXFILLER_103_0 vdd_d vss_d / DCAP64LVT
XXFILLER_103_64 vdd_d vss_d / DCAP64LVT
XXFILLER_103_128 vdd_d vss_d / DCAP64LVT
XXFILLER_103_192 vdd_d vss_d / DCAP64LVT
XXFILLER_103_256 vdd_d vss_d / DCAP64LVT
XXFILLER_103_320 vdd_d vss_d / DCAP64LVT
XXFILLER_103_384 vdd_d vss_d / DCAP64LVT
XXFILLER_103_448 vdd_d vss_d / DCAP64LVT
XXFILLER_103_512 vdd_d vss_d / DCAP64LVT
XXFILLER_103_576 vdd_d vss_d / DCAP64LVT
XXFILLER_103_640 vdd_d vss_d / DCAP64LVT
XXFILLER_103_704 vdd_d vss_d / DCAP64LVT
XXFILLER_103_768 vdd_d vss_d / DCAP64LVT
XXFILLER_103_832 vdd_d vss_d / DCAP64LVT
XXFILLER_103_896 vdd_d vss_d / DCAP64LVT
XXFILLER_103_960 vdd_d vss_d / DCAP64LVT
XXFILLER_103_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_103_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_103_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_103_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_103_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_103_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_103_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_103_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_103_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_103_1655 vdd_d vss_d / DCAP64LVT
XXFILLER_103_1788 vdd_d vss_d / DCAP64LVT
XXFILLER_103_1948 vdd_d vss_d / DCAP64LVT
XXFILLER_103_2012 vdd_d vss_d / DCAP64LVT
XXFILLER_103_2076 vdd_d vss_d / DCAP64LVT
XXFILLER_103_2140 vdd_d vss_d / DCAP64LVT
XXFILLER_103_2204 vdd_d vss_d / DCAP64LVT
XXFILLER_103_2268 vdd_d vss_d / DCAP64LVT
XXFILLER_104_0 vdd_d vss_d / DCAP64LVT
XXFILLER_104_64 vdd_d vss_d / DCAP64LVT
XXFILLER_104_128 vdd_d vss_d / DCAP64LVT
XXFILLER_104_192 vdd_d vss_d / DCAP64LVT
XXFILLER_104_256 vdd_d vss_d / DCAP64LVT
XXFILLER_104_320 vdd_d vss_d / DCAP64LVT
XXFILLER_104_384 vdd_d vss_d / DCAP64LVT
XXFILLER_104_448 vdd_d vss_d / DCAP64LVT
XXFILLER_104_512 vdd_d vss_d / DCAP64LVT
XXFILLER_104_576 vdd_d vss_d / DCAP64LVT
XXFILLER_104_640 vdd_d vss_d / DCAP64LVT
XXFILLER_104_704 vdd_d vss_d / DCAP64LVT
XXFILLER_104_768 vdd_d vss_d / DCAP64LVT
XXFILLER_104_832 vdd_d vss_d / DCAP64LVT
XXFILLER_104_896 vdd_d vss_d / DCAP64LVT
XXFILLER_104_960 vdd_d vss_d / DCAP64LVT
XXFILLER_104_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_104_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_104_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_104_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_104_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_104_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_104_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_104_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_104_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_104_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_104_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_104_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_104_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_104_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_104_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_104_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_104_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_104_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_104_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_104_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_105_0 vdd_d vss_d / DCAP64LVT
XXFILLER_105_64 vdd_d vss_d / DCAP64LVT
XXFILLER_105_128 vdd_d vss_d / DCAP64LVT
XXFILLER_105_192 vdd_d vss_d / DCAP64LVT
XXFILLER_105_256 vdd_d vss_d / DCAP64LVT
XXFILLER_105_320 vdd_d vss_d / DCAP64LVT
XXFILLER_105_384 vdd_d vss_d / DCAP64LVT
XXFILLER_105_448 vdd_d vss_d / DCAP64LVT
XXFILLER_105_512 vdd_d vss_d / DCAP64LVT
XXFILLER_105_576 vdd_d vss_d / DCAP64LVT
XXFILLER_105_640 vdd_d vss_d / DCAP64LVT
XXFILLER_105_704 vdd_d vss_d / DCAP64LVT
XXFILLER_105_768 vdd_d vss_d / DCAP64LVT
XXFILLER_105_832 vdd_d vss_d / DCAP64LVT
XXFILLER_105_896 vdd_d vss_d / DCAP64LVT
XXFILLER_105_960 vdd_d vss_d / DCAP64LVT
XXFILLER_105_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_105_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_105_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_105_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_105_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_105_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_105_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_105_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_105_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_105_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_105_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_105_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_105_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_105_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_105_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_105_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_105_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_105_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_105_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_105_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_106_0 vdd_d vss_d / DCAP64LVT
XXFILLER_106_64 vdd_d vss_d / DCAP64LVT
XXFILLER_106_128 vdd_d vss_d / DCAP64LVT
XXFILLER_106_192 vdd_d vss_d / DCAP64LVT
XXFILLER_106_256 vdd_d vss_d / DCAP64LVT
XXFILLER_106_320 vdd_d vss_d / DCAP64LVT
XXFILLER_106_384 vdd_d vss_d / DCAP64LVT
XXFILLER_106_448 vdd_d vss_d / DCAP64LVT
XXFILLER_106_512 vdd_d vss_d / DCAP64LVT
XXFILLER_106_576 vdd_d vss_d / DCAP64LVT
XXFILLER_106_640 vdd_d vss_d / DCAP64LVT
XXFILLER_106_704 vdd_d vss_d / DCAP64LVT
XXFILLER_106_768 vdd_d vss_d / DCAP64LVT
XXFILLER_106_832 vdd_d vss_d / DCAP64LVT
XXFILLER_106_896 vdd_d vss_d / DCAP64LVT
XXFILLER_106_960 vdd_d vss_d / DCAP64LVT
XXFILLER_106_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_106_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_106_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_106_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_106_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_106_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_106_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_106_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_106_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_106_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_106_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_106_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_106_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_106_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_106_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_106_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_106_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_106_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_106_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_106_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_107_0 vdd_d vss_d / DCAP64LVT
XXFILLER_107_64 vdd_d vss_d / DCAP64LVT
XXFILLER_107_128 vdd_d vss_d / DCAP64LVT
XXFILLER_107_192 vdd_d vss_d / DCAP64LVT
XXFILLER_107_256 vdd_d vss_d / DCAP64LVT
XXFILLER_107_320 vdd_d vss_d / DCAP64LVT
XXFILLER_107_384 vdd_d vss_d / DCAP64LVT
XXFILLER_107_448 vdd_d vss_d / DCAP64LVT
XXFILLER_107_512 vdd_d vss_d / DCAP64LVT
XXFILLER_107_576 vdd_d vss_d / DCAP64LVT
XXFILLER_107_640 vdd_d vss_d / DCAP64LVT
XXFILLER_107_704 vdd_d vss_d / DCAP64LVT
XXFILLER_107_768 vdd_d vss_d / DCAP64LVT
XXFILLER_107_832 vdd_d vss_d / DCAP64LVT
XXFILLER_107_896 vdd_d vss_d / DCAP64LVT
XXFILLER_107_960 vdd_d vss_d / DCAP64LVT
XXFILLER_107_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_107_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_107_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_107_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_107_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_107_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_107_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_107_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_107_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_107_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_107_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_107_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_107_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_107_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_107_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_107_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_107_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_107_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_107_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_107_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_108_0 vdd_d vss_d / DCAP64LVT
XXFILLER_108_64 vdd_d vss_d / DCAP64LVT
XXFILLER_108_128 vdd_d vss_d / DCAP64LVT
XXFILLER_108_192 vdd_d vss_d / DCAP64LVT
XXFILLER_108_256 vdd_d vss_d / DCAP64LVT
XXFILLER_108_320 vdd_d vss_d / DCAP64LVT
XXFILLER_108_384 vdd_d vss_d / DCAP64LVT
XXFILLER_108_448 vdd_d vss_d / DCAP64LVT
XXFILLER_108_512 vdd_d vss_d / DCAP64LVT
XXFILLER_108_576 vdd_d vss_d / DCAP64LVT
XXFILLER_108_640 vdd_d vss_d / DCAP64LVT
XXFILLER_108_704 vdd_d vss_d / DCAP64LVT
XXFILLER_108_768 vdd_d vss_d / DCAP64LVT
XXFILLER_108_832 vdd_d vss_d / DCAP64LVT
XXFILLER_108_942 vdd_d vss_d / DCAP64LVT
XXFILLER_108_1006 vdd_d vss_d / DCAP64LVT
XXFILLER_108_1070 vdd_d vss_d / DCAP64LVT
XXFILLER_108_1134 vdd_d vss_d / DCAP64LVT
XXFILLER_108_1198 vdd_d vss_d / DCAP64LVT
XXFILLER_108_1262 vdd_d vss_d / DCAP64LVT
XXFILLER_108_1326 vdd_d vss_d / DCAP64LVT
XXFILLER_108_1443 vdd_d vss_d / DCAP64LVT
XXFILLER_108_1507 vdd_d vss_d / DCAP64LVT
XXFILLER_108_1571 vdd_d vss_d / DCAP64LVT
XXFILLER_108_1635 vdd_d vss_d / DCAP64LVT
XXFILLER_108_1699 vdd_d vss_d / DCAP64LVT
XXFILLER_108_1763 vdd_d vss_d / DCAP64LVT
XXFILLER_108_1827 vdd_d vss_d / DCAP64LVT
XXFILLER_108_1891 vdd_d vss_d / DCAP64LVT
XXFILLER_108_1955 vdd_d vss_d / DCAP64LVT
XXFILLER_108_2019 vdd_d vss_d / DCAP64LVT
XXFILLER_108_2083 vdd_d vss_d / DCAP64LVT
XXFILLER_108_2147 vdd_d vss_d / DCAP64LVT
XXFILLER_108_2211 vdd_d vss_d / DCAP64LVT
XXFILLER_108_2275 vdd_d vss_d / DCAP64LVT
XXFILLER_109_0 vdd_d vss_d / DCAP64LVT
XXFILLER_109_64 vdd_d vss_d / DCAP64LVT
XXFILLER_109_128 vdd_d vss_d / DCAP64LVT
XXFILLER_109_192 vdd_d vss_d / DCAP64LVT
XXFILLER_109_256 vdd_d vss_d / DCAP64LVT
XXFILLER_109_320 vdd_d vss_d / DCAP64LVT
XXFILLER_109_384 vdd_d vss_d / DCAP64LVT
XXFILLER_109_448 vdd_d vss_d / DCAP64LVT
XXFILLER_109_512 vdd_d vss_d / DCAP64LVT
XXFILLER_109_576 vdd_d vss_d / DCAP64LVT
XXFILLER_109_640 vdd_d vss_d / DCAP64LVT
XXFILLER_109_704 vdd_d vss_d / DCAP64LVT
XXFILLER_109_768 vdd_d vss_d / DCAP64LVT
XXFILLER_109_832 vdd_d vss_d / DCAP64LVT
XXFILLER_109_896 vdd_d vss_d / DCAP64LVT
XXFILLER_109_960 vdd_d vss_d / DCAP64LVT
XXFILLER_109_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_109_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_109_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_109_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_109_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_109_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_109_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_109_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_109_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_109_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_109_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_109_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_109_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_109_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_109_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_109_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_109_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_109_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_109_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_109_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_110_0 vdd_d vss_d / DCAP64LVT
XXFILLER_110_64 vdd_d vss_d / DCAP64LVT
XXFILLER_110_128 vdd_d vss_d / DCAP64LVT
XXFILLER_110_192 vdd_d vss_d / DCAP64LVT
XXFILLER_110_256 vdd_d vss_d / DCAP64LVT
XXFILLER_110_320 vdd_d vss_d / DCAP64LVT
XXFILLER_110_384 vdd_d vss_d / DCAP64LVT
XXFILLER_110_448 vdd_d vss_d / DCAP64LVT
XXFILLER_110_512 vdd_d vss_d / DCAP64LVT
XXFILLER_110_576 vdd_d vss_d / DCAP64LVT
XXFILLER_110_640 vdd_d vss_d / DCAP64LVT
XXFILLER_110_704 vdd_d vss_d / DCAP64LVT
XXFILLER_110_768 vdd_d vss_d / DCAP64LVT
XXFILLER_110_832 vdd_d vss_d / DCAP64LVT
XXFILLER_110_896 vdd_d vss_d / DCAP64LVT
XXFILLER_110_960 vdd_d vss_d / DCAP64LVT
XXFILLER_110_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_110_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_110_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_110_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_110_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_110_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_110_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_110_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_110_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_110_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_110_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_110_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_110_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_110_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_110_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_110_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_110_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_110_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_110_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_110_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_111_0 vdd_d vss_d / DCAP64LVT
XXFILLER_111_64 vdd_d vss_d / DCAP64LVT
XXFILLER_111_128 vdd_d vss_d / DCAP64LVT
XXFILLER_111_192 vdd_d vss_d / DCAP64LVT
XXFILLER_111_256 vdd_d vss_d / DCAP64LVT
XXFILLER_111_320 vdd_d vss_d / DCAP64LVT
XXFILLER_111_384 vdd_d vss_d / DCAP64LVT
XXFILLER_111_448 vdd_d vss_d / DCAP64LVT
XXFILLER_111_512 vdd_d vss_d / DCAP64LVT
XXFILLER_111_576 vdd_d vss_d / DCAP64LVT
XXFILLER_111_640 vdd_d vss_d / DCAP64LVT
XXFILLER_111_704 vdd_d vss_d / DCAP64LVT
XXFILLER_111_768 vdd_d vss_d / DCAP64LVT
XXFILLER_111_832 vdd_d vss_d / DCAP64LVT
XXFILLER_111_919 vdd_d vss_d / DCAP64LVT
XXFILLER_111_983 vdd_d vss_d / DCAP64LVT
XXFILLER_111_1047 vdd_d vss_d / DCAP64LVT
XXFILLER_111_1111 vdd_d vss_d / DCAP64LVT
XXFILLER_111_1175 vdd_d vss_d / DCAP64LVT
XXFILLER_111_1239 vdd_d vss_d / DCAP64LVT
XXFILLER_111_1303 vdd_d vss_d / DCAP64LVT
XXFILLER_111_1367 vdd_d vss_d / DCAP64LVT
XXFILLER_111_1489 vdd_d vss_d / DCAP64LVT
XXFILLER_111_1553 vdd_d vss_d / DCAP64LVT
XXFILLER_111_1617 vdd_d vss_d / DCAP64LVT
XXFILLER_111_1681 vdd_d vss_d / DCAP64LVT
XXFILLER_111_1745 vdd_d vss_d / DCAP64LVT
XXFILLER_111_1901 vdd_d vss_d / DCAP64LVT
XXFILLER_111_1965 vdd_d vss_d / DCAP64LVT
XXFILLER_111_2029 vdd_d vss_d / DCAP64LVT
XXFILLER_111_2093 vdd_d vss_d / DCAP64LVT
XXFILLER_111_2157 vdd_d vss_d / DCAP64LVT
XXFILLER_111_2221 vdd_d vss_d / DCAP64LVT
XXFILLER_111_2285 vdd_d vss_d / DCAP64LVT
XXFILLER_112_0 vdd_d vss_d / DCAP64LVT
XXFILLER_112_64 vdd_d vss_d / DCAP64LVT
XXFILLER_112_128 vdd_d vss_d / DCAP64LVT
XXFILLER_112_192 vdd_d vss_d / DCAP64LVT
XXFILLER_112_587 vdd_d vss_d / DCAP64LVT
XXFILLER_112_651 vdd_d vss_d / DCAP64LVT
XXFILLER_112_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_112_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_112_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_112_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_112_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_112_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_112_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_112_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_113_0 vdd_d vss_d / DCAP64LVT
XXFILLER_113_64 vdd_d vss_d / DCAP64LVT
XXFILLER_113_128 vdd_d vss_d / DCAP64LVT
XXFILLER_113_192 vdd_d vss_d / DCAP64LVT
XXFILLER_113_587 vdd_d vss_d / DCAP64LVT
XXFILLER_113_651 vdd_d vss_d / DCAP64LVT
XXFILLER_113_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_113_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_113_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_113_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_113_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_113_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_113_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_113_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_114_0 vdd_d vss_d / DCAP64LVT
XXFILLER_114_64 vdd_d vss_d / DCAP64LVT
XXFILLER_114_128 vdd_d vss_d / DCAP64LVT
XXFILLER_114_192 vdd_d vss_d / DCAP64LVT
XXFILLER_114_587 vdd_d vss_d / DCAP64LVT
XXFILLER_114_651 vdd_d vss_d / DCAP64LVT
XXFILLER_114_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_114_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_114_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_114_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_114_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_114_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_114_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_114_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_115_0 vdd_d vss_d / DCAP64LVT
XXFILLER_115_64 vdd_d vss_d / DCAP64LVT
XXFILLER_115_128 vdd_d vss_d / DCAP64LVT
XXFILLER_115_192 vdd_d vss_d / DCAP64LVT
XXFILLER_115_587 vdd_d vss_d / DCAP64LVT
XXFILLER_115_651 vdd_d vss_d / DCAP64LVT
XXFILLER_115_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_115_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_115_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_115_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_115_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_115_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_115_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_115_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_116_0 vdd_d vss_d / DCAP64LVT
XXFILLER_116_64 vdd_d vss_d / DCAP64LVT
XXFILLER_116_128 vdd_d vss_d / DCAP64LVT
XXFILLER_116_192 vdd_d vss_d / DCAP64LVT
XXFILLER_116_587 vdd_d vss_d / DCAP64LVT
XXFILLER_116_651 vdd_d vss_d / DCAP64LVT
XXFILLER_116_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_116_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_116_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_116_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_116_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_116_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_116_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_116_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_117_0 vdd_d vss_d / DCAP64LVT
XXFILLER_117_64 vdd_d vss_d / DCAP64LVT
XXFILLER_117_128 vdd_d vss_d / DCAP64LVT
XXFILLER_117_192 vdd_d vss_d / DCAP64LVT
XXFILLER_117_587 vdd_d vss_d / DCAP64LVT
XXFILLER_117_651 vdd_d vss_d / DCAP64LVT
XXFILLER_117_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_117_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_117_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_117_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_117_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_117_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_117_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_117_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_118_0 vdd_d vss_d / DCAP64LVT
XXFILLER_118_64 vdd_d vss_d / DCAP64LVT
XXFILLER_118_128 vdd_d vss_d / DCAP64LVT
XXFILLER_118_192 vdd_d vss_d / DCAP64LVT
XXFILLER_118_587 vdd_d vss_d / DCAP64LVT
XXFILLER_118_651 vdd_d vss_d / DCAP64LVT
XXFILLER_118_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_118_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_118_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_118_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_118_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_118_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_118_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_118_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_119_0 vdd_d vss_d / DCAP64LVT
XXFILLER_119_64 vdd_d vss_d / DCAP64LVT
XXFILLER_119_128 vdd_d vss_d / DCAP64LVT
XXFILLER_119_192 vdd_d vss_d / DCAP64LVT
XXFILLER_119_587 vdd_d vss_d / DCAP64LVT
XXFILLER_119_651 vdd_d vss_d / DCAP64LVT
XXFILLER_119_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_119_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_119_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_119_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_119_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_119_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_119_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_119_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_120_0 vdd_d vss_d / DCAP64LVT
XXFILLER_120_64 vdd_d vss_d / DCAP64LVT
XXFILLER_120_128 vdd_d vss_d / DCAP64LVT
XXFILLER_120_192 vdd_d vss_d / DCAP64LVT
XXFILLER_120_587 vdd_d vss_d / DCAP64LVT
XXFILLER_120_651 vdd_d vss_d / DCAP64LVT
XXFILLER_120_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_120_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_120_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_120_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_120_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_120_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_120_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_120_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_121_0 vdd_d vss_d / DCAP64LVT
XXFILLER_121_64 vdd_d vss_d / DCAP64LVT
XXFILLER_121_128 vdd_d vss_d / DCAP64LVT
XXFILLER_121_192 vdd_d vss_d / DCAP64LVT
XXFILLER_121_587 vdd_d vss_d / DCAP64LVT
XXFILLER_121_651 vdd_d vss_d / DCAP64LVT
XXFILLER_121_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_121_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_121_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_121_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_121_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_121_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_121_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_121_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_122_0 vdd_d vss_d / DCAP64LVT
XXFILLER_122_64 vdd_d vss_d / DCAP64LVT
XXFILLER_122_128 vdd_d vss_d / DCAP64LVT
XXFILLER_122_192 vdd_d vss_d / DCAP64LVT
XXFILLER_122_587 vdd_d vss_d / DCAP64LVT
XXFILLER_122_651 vdd_d vss_d / DCAP64LVT
XXFILLER_122_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_122_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_122_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_122_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_122_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_122_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_122_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_122_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_123_0 vdd_d vss_d / DCAP64LVT
XXFILLER_123_64 vdd_d vss_d / DCAP64LVT
XXFILLER_123_128 vdd_d vss_d / DCAP64LVT
XXFILLER_123_192 vdd_d vss_d / DCAP64LVT
XXFILLER_123_587 vdd_d vss_d / DCAP64LVT
XXFILLER_123_651 vdd_d vss_d / DCAP64LVT
XXFILLER_123_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_123_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_123_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_123_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_123_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_123_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_123_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_123_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_124_0 vdd_d vss_d / DCAP64LVT
XXFILLER_124_64 vdd_d vss_d / DCAP64LVT
XXFILLER_124_128 vdd_d vss_d / DCAP64LVT
XXFILLER_124_192 vdd_d vss_d / DCAP64LVT
XXFILLER_124_587 vdd_d vss_d / DCAP64LVT
XXFILLER_124_651 vdd_d vss_d / DCAP64LVT
XXFILLER_124_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_124_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_124_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_124_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_124_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_124_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_124_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_124_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_125_0 vdd_d vss_d / DCAP64LVT
XXFILLER_125_64 vdd_d vss_d / DCAP64LVT
XXFILLER_125_128 vdd_d vss_d / DCAP64LVT
XXFILLER_125_192 vdd_d vss_d / DCAP64LVT
XXFILLER_125_587 vdd_d vss_d / DCAP64LVT
XXFILLER_125_651 vdd_d vss_d / DCAP64LVT
XXFILLER_125_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_125_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_125_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_125_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_125_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_125_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_125_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_125_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_126_0 vdd_d vss_d / DCAP64LVT
XXFILLER_126_64 vdd_d vss_d / DCAP64LVT
XXFILLER_126_128 vdd_d vss_d / DCAP64LVT
XXFILLER_126_192 vdd_d vss_d / DCAP64LVT
XXFILLER_126_587 vdd_d vss_d / DCAP64LVT
XXFILLER_126_651 vdd_d vss_d / DCAP64LVT
XXFILLER_126_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_126_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_126_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_126_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_126_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_126_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_126_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_126_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_127_0 vdd_d vss_d / DCAP64LVT
XXFILLER_127_64 vdd_d vss_d / DCAP64LVT
XXFILLER_127_128 vdd_d vss_d / DCAP64LVT
XXFILLER_127_192 vdd_d vss_d / DCAP64LVT
XXFILLER_127_587 vdd_d vss_d / DCAP64LVT
XXFILLER_127_651 vdd_d vss_d / DCAP64LVT
XXFILLER_127_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_127_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_127_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_127_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_127_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_127_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_127_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_127_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_128_0 vdd_d vss_d / DCAP64LVT
XXFILLER_128_64 vdd_d vss_d / DCAP64LVT
XXFILLER_128_128 vdd_d vss_d / DCAP64LVT
XXFILLER_128_192 vdd_d vss_d / DCAP64LVT
XXFILLER_128_587 vdd_d vss_d / DCAP64LVT
XXFILLER_128_651 vdd_d vss_d / DCAP64LVT
XXFILLER_128_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_128_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_128_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_128_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_128_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_128_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_128_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_128_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_129_0 vdd_d vss_d / DCAP64LVT
XXFILLER_129_64 vdd_d vss_d / DCAP64LVT
XXFILLER_129_128 vdd_d vss_d / DCAP64LVT
XXFILLER_129_192 vdd_d vss_d / DCAP64LVT
XXFILLER_129_587 vdd_d vss_d / DCAP64LVT
XXFILLER_129_651 vdd_d vss_d / DCAP64LVT
XXFILLER_129_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_129_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_129_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_129_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_129_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_129_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_129_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_129_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_130_0 vdd_d vss_d / DCAP64LVT
XXFILLER_130_64 vdd_d vss_d / DCAP64LVT
XXFILLER_130_128 vdd_d vss_d / DCAP64LVT
XXFILLER_130_192 vdd_d vss_d / DCAP64LVT
XXFILLER_130_587 vdd_d vss_d / DCAP64LVT
XXFILLER_130_651 vdd_d vss_d / DCAP64LVT
XXFILLER_130_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_130_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_130_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_130_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_130_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_130_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_130_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_130_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_131_0 vdd_d vss_d / DCAP64LVT
XXFILLER_131_64 vdd_d vss_d / DCAP64LVT
XXFILLER_131_128 vdd_d vss_d / DCAP64LVT
XXFILLER_131_587 vdd_d vss_d / DCAP64LVT
XXFILLER_131_651 vdd_d vss_d / DCAP64LVT
XXFILLER_131_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_131_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_131_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_131_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_131_2099 vdd_d vss_d / DCAP64LVT
XXFILLER_131_2163 vdd_d vss_d / DCAP64LVT
XXFILLER_131_2227 vdd_d vss_d / DCAP64LVT
XXFILLER_132_0 vdd_d vss_d / DCAP64LVT
XXFILLER_132_64 vdd_d vss_d / DCAP64LVT
XXFILLER_132_128 vdd_d vss_d / DCAP64LVT
XXFILLER_132_192 vdd_d vss_d / DCAP64LVT
XXFILLER_132_587 vdd_d vss_d / DCAP64LVT
XXFILLER_132_651 vdd_d vss_d / DCAP64LVT
XXFILLER_132_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_132_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_132_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_132_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_132_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_132_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_132_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_132_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_133_0 vdd_d vss_d / DCAP64LVT
XXFILLER_133_64 vdd_d vss_d / DCAP64LVT
XXFILLER_133_128 vdd_d vss_d / DCAP64LVT
XXFILLER_133_192 vdd_d vss_d / DCAP64LVT
XXFILLER_133_587 vdd_d vss_d / DCAP64LVT
XXFILLER_133_651 vdd_d vss_d / DCAP64LVT
XXFILLER_133_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_133_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_133_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_133_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_133_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_133_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_133_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_133_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_134_0 vdd_d vss_d / DCAP64LVT
XXFILLER_134_64 vdd_d vss_d / DCAP64LVT
XXFILLER_134_128 vdd_d vss_d / DCAP64LVT
XXFILLER_134_192 vdd_d vss_d / DCAP64LVT
XXFILLER_134_587 vdd_d vss_d / DCAP64LVT
XXFILLER_134_651 vdd_d vss_d / DCAP64LVT
XXFILLER_134_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_134_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_134_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_134_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_134_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_134_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_134_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_134_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_135_0 vdd_d vss_d / DCAP64LVT
XXFILLER_135_64 vdd_d vss_d / DCAP64LVT
XXFILLER_135_128 vdd_d vss_d / DCAP64LVT
XXFILLER_135_192 vdd_d vss_d / DCAP64LVT
XXFILLER_135_587 vdd_d vss_d / DCAP64LVT
XXFILLER_135_651 vdd_d vss_d / DCAP64LVT
XXFILLER_135_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_135_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_135_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_135_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_135_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_135_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_135_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_135_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_136_0 vdd_d vss_d / DCAP64LVT
XXFILLER_136_64 vdd_d vss_d / DCAP64LVT
XXFILLER_136_128 vdd_d vss_d / DCAP64LVT
XXFILLER_136_192 vdd_d vss_d / DCAP64LVT
XXFILLER_136_587 vdd_d vss_d / DCAP64LVT
XXFILLER_136_651 vdd_d vss_d / DCAP64LVT
XXFILLER_136_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_136_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_136_1637 vdd_d vss_d / DCAP64LVT
XXFILLER_136_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_136_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_136_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_136_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_137_0 vdd_d vss_d / DCAP64LVT
XXFILLER_137_64 vdd_d vss_d / DCAP64LVT
XXFILLER_137_128 vdd_d vss_d / DCAP64LVT
XXFILLER_137_192 vdd_d vss_d / DCAP64LVT
XXFILLER_137_587 vdd_d vss_d / DCAP64LVT
XXFILLER_137_651 vdd_d vss_d / DCAP64LVT
XXFILLER_137_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_137_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_137_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_137_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_137_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_137_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_137_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_137_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_138_0 vdd_d vss_d / DCAP64LVT
XXFILLER_138_64 vdd_d vss_d / DCAP64LVT
XXFILLER_138_128 vdd_d vss_d / DCAP64LVT
XXFILLER_138_192 vdd_d vss_d / DCAP64LVT
XXFILLER_138_587 vdd_d vss_d / DCAP64LVT
XXFILLER_138_651 vdd_d vss_d / DCAP64LVT
XXFILLER_138_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_138_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_138_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_138_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_138_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_138_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_138_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_138_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_139_0 vdd_d vss_d / DCAP64LVT
XXFILLER_139_64 vdd_d vss_d / DCAP64LVT
XXFILLER_139_128 vdd_d vss_d / DCAP64LVT
XXFILLER_139_192 vdd_d vss_d / DCAP64LVT
XXFILLER_139_587 vdd_d vss_d / DCAP64LVT
XXFILLER_139_651 vdd_d vss_d / DCAP64LVT
XXFILLER_139_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_139_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_139_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_139_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_139_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_139_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_139_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_139_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_140_0 vdd_d vss_d / DCAP64LVT
XXFILLER_140_64 vdd_d vss_d / DCAP64LVT
XXFILLER_140_128 vdd_d vss_d / DCAP64LVT
XXFILLER_140_192 vdd_d vss_d / DCAP64LVT
XXFILLER_140_587 vdd_d vss_d / DCAP64LVT
XXFILLER_140_651 vdd_d vss_d / DCAP64LVT
XXFILLER_140_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_140_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_140_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_140_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_140_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_140_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_140_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_141_0 vdd_d vss_d / DCAP64LVT
XXFILLER_141_64 vdd_d vss_d / DCAP64LVT
XXFILLER_141_128 vdd_d vss_d / DCAP64LVT
XXFILLER_141_192 vdd_d vss_d / DCAP64LVT
XXFILLER_141_587 vdd_d vss_d / DCAP64LVT
XXFILLER_141_651 vdd_d vss_d / DCAP64LVT
XXFILLER_141_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_141_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_141_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_141_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_141_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_141_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_141_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_142_0 vdd_d vss_d / DCAP64LVT
XXFILLER_142_64 vdd_d vss_d / DCAP64LVT
XXFILLER_142_128 vdd_d vss_d / DCAP64LVT
XXFILLER_142_192 vdd_d vss_d / DCAP64LVT
XXFILLER_142_587 vdd_d vss_d / DCAP64LVT
XXFILLER_142_651 vdd_d vss_d / DCAP64LVT
XXFILLER_142_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_142_1199 vdd_d vss_d / DCAP64LVT
XXFILLER_142_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_142_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_142_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_142_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_142_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_142_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_143_0 vdd_d vss_d / DCAP64LVT
XXFILLER_143_64 vdd_d vss_d / DCAP64LVT
XXFILLER_143_128 vdd_d vss_d / DCAP64LVT
XXFILLER_143_192 vdd_d vss_d / DCAP64LVT
XXFILLER_143_587 vdd_d vss_d / DCAP64LVT
XXFILLER_143_651 vdd_d vss_d / DCAP64LVT
XXFILLER_143_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_143_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_143_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_143_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_143_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_143_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_143_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_143_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_144_0 vdd_d vss_d / DCAP64LVT
XXFILLER_144_64 vdd_d vss_d / DCAP64LVT
XXFILLER_144_128 vdd_d vss_d / DCAP64LVT
XXFILLER_144_192 vdd_d vss_d / DCAP64LVT
XXFILLER_144_587 vdd_d vss_d / DCAP64LVT
XXFILLER_144_651 vdd_d vss_d / DCAP64LVT
XXFILLER_144_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_144_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_144_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_144_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_144_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_144_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_144_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_144_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_145_0 vdd_d vss_d / DCAP64LVT
XXFILLER_145_64 vdd_d vss_d / DCAP64LVT
XXFILLER_145_128 vdd_d vss_d / DCAP64LVT
XXFILLER_145_192 vdd_d vss_d / DCAP64LVT
XXFILLER_145_587 vdd_d vss_d / DCAP64LVT
XXFILLER_145_651 vdd_d vss_d / DCAP64LVT
XXFILLER_145_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_145_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_145_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_145_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_145_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_145_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_145_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_145_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_146_0 vdd_d vss_d / DCAP64LVT
XXFILLER_146_64 vdd_d vss_d / DCAP64LVT
XXFILLER_146_128 vdd_d vss_d / DCAP64LVT
XXFILLER_146_192 vdd_d vss_d / DCAP64LVT
XXFILLER_146_587 vdd_d vss_d / DCAP64LVT
XXFILLER_146_651 vdd_d vss_d / DCAP64LVT
XXFILLER_146_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_146_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_146_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_146_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_146_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_146_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_146_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_146_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_147_0 vdd_d vss_d / DCAP64LVT
XXFILLER_147_64 vdd_d vss_d / DCAP64LVT
XXFILLER_147_128 vdd_d vss_d / DCAP64LVT
XXFILLER_147_192 vdd_d vss_d / DCAP64LVT
XXFILLER_147_587 vdd_d vss_d / DCAP64LVT
XXFILLER_147_651 vdd_d vss_d / DCAP64LVT
XXFILLER_147_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_147_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_147_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_147_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_147_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_147_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_147_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_147_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_148_0 vdd_d vss_d / DCAP64LVT
XXFILLER_148_64 vdd_d vss_d / DCAP64LVT
XXFILLER_148_128 vdd_d vss_d / DCAP64LVT
XXFILLER_148_192 vdd_d vss_d / DCAP64LVT
XXFILLER_148_587 vdd_d vss_d / DCAP64LVT
XXFILLER_148_651 vdd_d vss_d / DCAP64LVT
XXFILLER_148_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_148_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_148_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_148_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_148_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_148_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_148_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_148_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_149_0 vdd_d vss_d / DCAP64LVT
XXFILLER_149_64 vdd_d vss_d / DCAP64LVT
XXFILLER_149_128 vdd_d vss_d / DCAP64LVT
XXFILLER_149_192 vdd_d vss_d / DCAP64LVT
XXFILLER_149_587 vdd_d vss_d / DCAP64LVT
XXFILLER_149_651 vdd_d vss_d / DCAP64LVT
XXFILLER_149_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_149_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_149_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_149_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_149_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_149_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_149_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_149_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_150_0 vdd_d vss_d / DCAP64LVT
XXFILLER_150_64 vdd_d vss_d / DCAP64LVT
XXFILLER_150_128 vdd_d vss_d / DCAP64LVT
XXFILLER_150_192 vdd_d vss_d / DCAP64LVT
XXFILLER_150_256 vdd_d vss_d / DCAP64LVT
XXFILLER_150_320 vdd_d vss_d / DCAP64LVT
XXFILLER_150_448 vdd_d vss_d / DCAP64LVT
XXFILLER_150_512 vdd_d vss_d / DCAP64LVT
XXFILLER_150_576 vdd_d vss_d / DCAP64LVT
XXFILLER_150_640 vdd_d vss_d / DCAP64LVT
XXFILLER_150_704 vdd_d vss_d / DCAP64LVT
XXFILLER_150_768 vdd_d vss_d / DCAP64LVT
XXFILLER_150_832 vdd_d vss_d / DCAP64LVT
XXFILLER_150_896 vdd_d vss_d / DCAP64LVT
XXFILLER_150_960 vdd_d vss_d / DCAP64LVT
XXFILLER_150_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_150_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_150_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_150_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_150_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_150_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_150_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_150_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_150_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_150_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_150_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_150_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_150_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_150_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_150_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_150_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_150_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_150_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_150_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_150_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_151_0 vdd_d vss_d / DCAP64LVT
XXFILLER_151_64 vdd_d vss_d / DCAP64LVT
XXFILLER_151_128 vdd_d vss_d / DCAP64LVT
XXFILLER_151_192 vdd_d vss_d / DCAP64LVT
XXFILLER_151_256 vdd_d vss_d / DCAP64LVT
XXFILLER_151_320 vdd_d vss_d / DCAP64LVT
XXFILLER_151_456 vdd_d vss_d / DCAP64LVT
XXFILLER_151_520 vdd_d vss_d / DCAP64LVT
XXFILLER_151_584 vdd_d vss_d / DCAP64LVT
XXFILLER_151_648 vdd_d vss_d / DCAP64LVT
XXFILLER_151_712 vdd_d vss_d / DCAP64LVT
XXFILLER_151_776 vdd_d vss_d / DCAP64LVT
XXFILLER_151_840 vdd_d vss_d / DCAP64LVT
XXFILLER_151_975 vdd_d vss_d / DCAP64LVT
XXFILLER_151_1039 vdd_d vss_d / DCAP64LVT
XXFILLER_151_1103 vdd_d vss_d / DCAP64LVT
XXFILLER_151_1167 vdd_d vss_d / DCAP64LVT
XXFILLER_151_1231 vdd_d vss_d / DCAP64LVT
XXFILLER_151_1295 vdd_d vss_d / DCAP64LVT
XXFILLER_151_1443 vdd_d vss_d / DCAP64LVT
XXFILLER_151_1507 vdd_d vss_d / DCAP64LVT
XXFILLER_151_1571 vdd_d vss_d / DCAP64LVT
XXFILLER_151_1635 vdd_d vss_d / DCAP64LVT
XXFILLER_151_1699 vdd_d vss_d / DCAP64LVT
XXFILLER_151_1763 vdd_d vss_d / DCAP64LVT
XXFILLER_151_1827 vdd_d vss_d / DCAP64LVT
XXFILLER_151_1934 vdd_d vss_d / DCAP64LVT
XXFILLER_151_1998 vdd_d vss_d / DCAP64LVT
XXFILLER_151_2062 vdd_d vss_d / DCAP64LVT
XXFILLER_151_2126 vdd_d vss_d / DCAP64LVT
XXFILLER_151_2190 vdd_d vss_d / DCAP64LVT
XXFILLER_151_2254 vdd_d vss_d / DCAP64LVT
XXFILLER_152_0 vdd_d vss_d / DCAP64LVT
XXFILLER_152_64 vdd_d vss_d / DCAP64LVT
XXFILLER_152_128 vdd_d vss_d / DCAP64LVT
XXFILLER_152_192 vdd_d vss_d / DCAP64LVT
XXFILLER_152_256 vdd_d vss_d / DCAP64LVT
XXFILLER_152_320 vdd_d vss_d / DCAP64LVT
XXFILLER_152_384 vdd_d vss_d / DCAP64LVT
XXFILLER_152_448 vdd_d vss_d / DCAP64LVT
XXFILLER_152_512 vdd_d vss_d / DCAP64LVT
XXFILLER_152_576 vdd_d vss_d / DCAP64LVT
XXFILLER_152_640 vdd_d vss_d / DCAP64LVT
XXFILLER_152_704 vdd_d vss_d / DCAP64LVT
XXFILLER_152_768 vdd_d vss_d / DCAP64LVT
XXFILLER_152_832 vdd_d vss_d / DCAP64LVT
XXFILLER_152_896 vdd_d vss_d / DCAP64LVT
XXFILLER_152_960 vdd_d vss_d / DCAP64LVT
XXFILLER_152_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_152_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_152_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_152_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_152_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_152_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_152_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_152_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_152_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_152_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_152_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_152_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_152_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_152_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_152_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_152_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_152_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_152_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_152_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_152_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_153_0 vdd_d vss_d / DCAP64LVT
XXFILLER_153_64 vdd_d vss_d / DCAP64LVT
XXFILLER_153_128 vdd_d vss_d / DCAP64LVT
XXFILLER_153_192 vdd_d vss_d / DCAP64LVT
XXFILLER_153_256 vdd_d vss_d / DCAP64LVT
XXFILLER_153_320 vdd_d vss_d / DCAP64LVT
XXFILLER_153_384 vdd_d vss_d / DCAP64LVT
XXFILLER_153_448 vdd_d vss_d / DCAP64LVT
XXFILLER_153_512 vdd_d vss_d / DCAP64LVT
XXFILLER_153_576 vdd_d vss_d / DCAP64LVT
XXFILLER_153_640 vdd_d vss_d / DCAP64LVT
XXFILLER_153_704 vdd_d vss_d / DCAP64LVT
XXFILLER_153_768 vdd_d vss_d / DCAP64LVT
XXFILLER_153_832 vdd_d vss_d / DCAP64LVT
XXFILLER_153_896 vdd_d vss_d / DCAP64LVT
XXFILLER_153_960 vdd_d vss_d / DCAP64LVT
XXFILLER_153_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_153_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_153_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_153_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_153_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_153_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_153_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_153_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_153_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_153_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_153_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_153_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_153_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_153_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_153_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_153_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_153_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_153_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_153_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_153_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_154_0 vdd_d vss_d / DCAP64LVT
XXFILLER_154_64 vdd_d vss_d / DCAP64LVT
XXFILLER_154_128 vdd_d vss_d / DCAP64LVT
XXFILLER_154_192 vdd_d vss_d / DCAP64LVT
XXFILLER_154_256 vdd_d vss_d / DCAP64LVT
XXFILLER_154_320 vdd_d vss_d / DCAP64LVT
XXFILLER_154_384 vdd_d vss_d / DCAP64LVT
XXFILLER_154_448 vdd_d vss_d / DCAP64LVT
XXFILLER_154_512 vdd_d vss_d / DCAP64LVT
XXFILLER_154_576 vdd_d vss_d / DCAP64LVT
XXFILLER_154_640 vdd_d vss_d / DCAP64LVT
XXFILLER_154_704 vdd_d vss_d / DCAP64LVT
XXFILLER_154_768 vdd_d vss_d / DCAP64LVT
XXFILLER_154_832 vdd_d vss_d / DCAP64LVT
XXFILLER_154_896 vdd_d vss_d / DCAP64LVT
XXFILLER_154_960 vdd_d vss_d / DCAP64LVT
XXFILLER_154_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_154_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_154_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_154_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_154_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_154_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_154_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_154_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_154_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_154_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_154_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_154_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_154_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_154_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_154_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_154_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_154_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_154_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_154_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_154_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_155_0 vdd_d vss_d / DCAP64LVT
XXFILLER_155_64 vdd_d vss_d / DCAP64LVT
XXFILLER_155_128 vdd_d vss_d / DCAP64LVT
XXFILLER_155_192 vdd_d vss_d / DCAP64LVT
XXFILLER_155_256 vdd_d vss_d / DCAP64LVT
XXFILLER_155_320 vdd_d vss_d / DCAP64LVT
XXFILLER_155_384 vdd_d vss_d / DCAP64LVT
XXFILLER_155_448 vdd_d vss_d / DCAP64LVT
XXFILLER_155_512 vdd_d vss_d / DCAP64LVT
XXFILLER_155_576 vdd_d vss_d / DCAP64LVT
XXFILLER_155_640 vdd_d vss_d / DCAP64LVT
XXFILLER_155_704 vdd_d vss_d / DCAP64LVT
XXFILLER_155_768 vdd_d vss_d / DCAP64LVT
XXFILLER_155_832 vdd_d vss_d / DCAP64LVT
XXFILLER_155_896 vdd_d vss_d / DCAP64LVT
XXFILLER_155_960 vdd_d vss_d / DCAP64LVT
XXFILLER_155_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_155_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_155_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_155_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_155_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_155_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_155_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_155_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_155_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_155_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_155_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_155_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_155_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_155_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_155_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_155_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_155_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_155_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_155_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_155_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_156_0 vdd_d vss_d / DCAP64LVT
XXFILLER_156_64 vdd_d vss_d / DCAP64LVT
XXFILLER_156_128 vdd_d vss_d / DCAP64LVT
XXFILLER_156_192 vdd_d vss_d / DCAP64LVT
XXFILLER_156_256 vdd_d vss_d / DCAP64LVT
XXFILLER_156_320 vdd_d vss_d / DCAP64LVT
XXFILLER_156_384 vdd_d vss_d / DCAP64LVT
XXFILLER_156_448 vdd_d vss_d / DCAP64LVT
XXFILLER_156_512 vdd_d vss_d / DCAP64LVT
XXFILLER_156_576 vdd_d vss_d / DCAP64LVT
XXFILLER_156_640 vdd_d vss_d / DCAP64LVT
XXFILLER_156_704 vdd_d vss_d / DCAP64LVT
XXFILLER_156_768 vdd_d vss_d / DCAP64LVT
XXFILLER_156_832 vdd_d vss_d / DCAP64LVT
XXFILLER_156_896 vdd_d vss_d / DCAP64LVT
XXFILLER_156_960 vdd_d vss_d / DCAP64LVT
XXFILLER_156_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_156_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_156_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_156_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_156_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_156_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_156_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_156_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_156_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_156_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_156_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_156_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_156_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_156_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_156_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_156_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_156_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_156_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_156_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_156_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_157_0 vdd_d vss_d / DCAP64LVT
XXFILLER_157_64 vdd_d vss_d / DCAP64LVT
XXFILLER_157_128 vdd_d vss_d / DCAP64LVT
XXFILLER_157_192 vdd_d vss_d / DCAP64LVT
XXFILLER_157_256 vdd_d vss_d / DCAP64LVT
XXFILLER_157_320 vdd_d vss_d / DCAP64LVT
XXFILLER_157_384 vdd_d vss_d / DCAP64LVT
XXFILLER_157_448 vdd_d vss_d / DCAP64LVT
XXFILLER_157_512 vdd_d vss_d / DCAP64LVT
XXFILLER_157_576 vdd_d vss_d / DCAP64LVT
XXFILLER_157_640 vdd_d vss_d / DCAP64LVT
XXFILLER_157_704 vdd_d vss_d / DCAP64LVT
XXFILLER_157_768 vdd_d vss_d / DCAP64LVT
XXFILLER_157_832 vdd_d vss_d / DCAP64LVT
XXFILLER_157_896 vdd_d vss_d / DCAP64LVT
XXFILLER_157_960 vdd_d vss_d / DCAP64LVT
XXFILLER_157_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_157_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_157_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_157_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_157_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_157_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_157_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_157_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_157_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_157_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_157_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_157_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_157_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_157_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_157_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_157_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_157_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_157_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_157_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_157_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_158_0 vdd_d vss_d / DCAP64LVT
XXFILLER_158_64 vdd_d vss_d / DCAP64LVT
XXFILLER_158_128 vdd_d vss_d / DCAP64LVT
XXFILLER_158_192 vdd_d vss_d / DCAP64LVT
XXFILLER_158_256 vdd_d vss_d / DCAP64LVT
XXFILLER_158_320 vdd_d vss_d / DCAP64LVT
XXFILLER_158_384 vdd_d vss_d / DCAP64LVT
XXFILLER_158_448 vdd_d vss_d / DCAP64LVT
XXFILLER_158_512 vdd_d vss_d / DCAP64LVT
XXFILLER_158_576 vdd_d vss_d / DCAP64LVT
XXFILLER_158_706 vdd_d vss_d / DCAP64LVT
XXFILLER_158_770 vdd_d vss_d / DCAP64LVT
XXFILLER_158_834 vdd_d vss_d / DCAP64LVT
XXFILLER_158_898 vdd_d vss_d / DCAP64LVT
XXFILLER_158_962 vdd_d vss_d / DCAP64LVT
XXFILLER_158_1026 vdd_d vss_d / DCAP64LVT
XXFILLER_158_1090 vdd_d vss_d / DCAP64LVT
XXFILLER_158_1154 vdd_d vss_d / DCAP64LVT
XXFILLER_158_1218 vdd_d vss_d / DCAP64LVT
XXFILLER_158_1282 vdd_d vss_d / DCAP64LVT
XXFILLER_158_1346 vdd_d vss_d / DCAP64LVT
XXFILLER_158_1410 vdd_d vss_d / DCAP64LVT
XXFILLER_158_1474 vdd_d vss_d / DCAP64LVT
XXFILLER_158_1538 vdd_d vss_d / DCAP64LVT
XXFILLER_158_1602 vdd_d vss_d / DCAP64LVT
XXFILLER_158_1666 vdd_d vss_d / DCAP64LVT
XXFILLER_158_1730 vdd_d vss_d / DCAP64LVT
XXFILLER_158_1794 vdd_d vss_d / DCAP64LVT
XXFILLER_158_1858 vdd_d vss_d / DCAP64LVT
XXFILLER_158_1922 vdd_d vss_d / DCAP64LVT
XXFILLER_158_1986 vdd_d vss_d / DCAP64LVT
XXFILLER_158_2050 vdd_d vss_d / DCAP64LVT
XXFILLER_158_2114 vdd_d vss_d / DCAP64LVT
XXFILLER_158_2178 vdd_d vss_d / DCAP64LVT
XXFILLER_158_2242 vdd_d vss_d / DCAP64LVT
XXFILLER_159_0 vdd_d vss_d / DCAP64LVT
XXFILLER_159_64 vdd_d vss_d / DCAP64LVT
XXFILLER_159_128 vdd_d vss_d / DCAP64LVT
XXFILLER_159_192 vdd_d vss_d / DCAP64LVT
XXFILLER_159_256 vdd_d vss_d / DCAP64LVT
XXFILLER_159_320 vdd_d vss_d / DCAP64LVT
XXFILLER_159_384 vdd_d vss_d / DCAP64LVT
XXFILLER_159_448 vdd_d vss_d / DCAP64LVT
XXFILLER_159_512 vdd_d vss_d / DCAP64LVT
XXFILLER_159_576 vdd_d vss_d / DCAP64LVT
XXFILLER_159_640 vdd_d vss_d / DCAP64LVT
XXFILLER_159_704 vdd_d vss_d / DCAP64LVT
XXFILLER_159_768 vdd_d vss_d / DCAP64LVT
XXFILLER_159_832 vdd_d vss_d / DCAP64LVT
XXFILLER_159_896 vdd_d vss_d / DCAP64LVT
XXFILLER_159_960 vdd_d vss_d / DCAP64LVT
XXFILLER_159_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_159_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_159_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_159_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_159_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_159_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_159_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_159_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_159_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_159_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_159_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_159_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_159_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_159_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_159_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_159_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_159_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_159_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_159_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_159_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_160_0 vdd_d vss_d / DCAP64LVT
XXFILLER_160_64 vdd_d vss_d / DCAP64LVT
XXFILLER_160_128 vdd_d vss_d / DCAP64LVT
XXFILLER_160_192 vdd_d vss_d / DCAP64LVT
XXFILLER_160_256 vdd_d vss_d / DCAP64LVT
XXFILLER_160_320 vdd_d vss_d / DCAP64LVT
XXFILLER_160_384 vdd_d vss_d / DCAP64LVT
XXFILLER_160_448 vdd_d vss_d / DCAP64LVT
XXFILLER_160_512 vdd_d vss_d / DCAP64LVT
XXFILLER_160_576 vdd_d vss_d / DCAP64LVT
XXFILLER_160_640 vdd_d vss_d / DCAP64LVT
XXFILLER_160_704 vdd_d vss_d / DCAP64LVT
XXFILLER_160_768 vdd_d vss_d / DCAP64LVT
XXFILLER_160_832 vdd_d vss_d / DCAP64LVT
XXFILLER_160_896 vdd_d vss_d / DCAP64LVT
XXFILLER_160_960 vdd_d vss_d / DCAP64LVT
XXFILLER_160_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_160_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_160_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_160_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_160_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_160_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_160_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_160_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_160_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_160_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_160_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_160_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_160_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_160_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_160_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_160_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_160_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_160_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_160_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_160_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_161_0 vdd_d vss_d / DCAP64LVT
XXFILLER_161_64 vdd_d vss_d / DCAP64LVT
XXFILLER_161_128 vdd_d vss_d / DCAP64LVT
XXFILLER_161_192 vdd_d vss_d / DCAP64LVT
XXFILLER_161_256 vdd_d vss_d / DCAP64LVT
XXFILLER_161_320 vdd_d vss_d / DCAP64LVT
XXFILLER_161_384 vdd_d vss_d / DCAP64LVT
XXFILLER_161_448 vdd_d vss_d / DCAP64LVT
XXFILLER_161_512 vdd_d vss_d / DCAP64LVT
XXFILLER_161_576 vdd_d vss_d / DCAP64LVT
XXFILLER_161_640 vdd_d vss_d / DCAP64LVT
XXFILLER_161_704 vdd_d vss_d / DCAP64LVT
XXFILLER_161_768 vdd_d vss_d / DCAP64LVT
XXFILLER_161_832 vdd_d vss_d / DCAP64LVT
XXFILLER_161_896 vdd_d vss_d / DCAP64LVT
XXFILLER_161_960 vdd_d vss_d / DCAP64LVT
XXFILLER_161_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_161_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_161_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_161_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_161_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_161_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_161_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_161_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_161_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_161_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_161_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_161_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_161_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_161_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_161_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_161_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_161_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_161_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_161_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_161_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_162_0 vdd_d vss_d / DCAP64LVT
XXFILLER_162_64 vdd_d vss_d / DCAP64LVT
XXFILLER_162_128 vdd_d vss_d / DCAP64LVT
XXFILLER_162_192 vdd_d vss_d / DCAP64LVT
XXFILLER_162_256 vdd_d vss_d / DCAP64LVT
XXFILLER_162_320 vdd_d vss_d / DCAP64LVT
XXFILLER_162_384 vdd_d vss_d / DCAP64LVT
XXFILLER_162_448 vdd_d vss_d / DCAP64LVT
XXFILLER_162_512 vdd_d vss_d / DCAP64LVT
XXFILLER_162_576 vdd_d vss_d / DCAP64LVT
XXFILLER_162_640 vdd_d vss_d / DCAP64LVT
XXFILLER_162_704 vdd_d vss_d / DCAP64LVT
XXFILLER_162_768 vdd_d vss_d / DCAP64LVT
XXFILLER_162_832 vdd_d vss_d / DCAP64LVT
XXFILLER_162_896 vdd_d vss_d / DCAP64LVT
XXFILLER_162_960 vdd_d vss_d / DCAP64LVT
XXFILLER_162_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_162_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_162_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_162_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_162_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_162_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_162_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_162_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_162_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_162_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_162_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_162_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_162_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_162_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_162_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_162_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_162_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_162_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_162_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_162_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_163_0 vdd_d vss_d / DCAP64LVT
XXFILLER_163_64 vdd_d vss_d / DCAP64LVT
XXFILLER_163_128 vdd_d vss_d / DCAP64LVT
XXFILLER_163_192 vdd_d vss_d / DCAP64LVT
XXFILLER_163_256 vdd_d vss_d / DCAP64LVT
XXFILLER_163_320 vdd_d vss_d / DCAP64LVT
XXFILLER_163_384 vdd_d vss_d / DCAP64LVT
XXFILLER_163_448 vdd_d vss_d / DCAP64LVT
XXFILLER_163_512 vdd_d vss_d / DCAP64LVT
XXFILLER_163_576 vdd_d vss_d / DCAP64LVT
XXFILLER_163_640 vdd_d vss_d / DCAP64LVT
XXFILLER_163_704 vdd_d vss_d / DCAP64LVT
XXFILLER_163_768 vdd_d vss_d / DCAP64LVT
XXFILLER_163_832 vdd_d vss_d / DCAP64LVT
XXFILLER_163_896 vdd_d vss_d / DCAP64LVT
XXFILLER_163_960 vdd_d vss_d / DCAP64LVT
XXFILLER_163_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_163_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_163_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_163_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_163_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_163_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_163_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_163_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_163_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_163_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_163_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_163_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_163_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_163_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_163_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_163_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_163_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_163_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_163_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_163_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_164_0 vdd_d vss_d / DCAP64LVT
XXFILLER_164_64 vdd_d vss_d / DCAP64LVT
XXFILLER_164_128 vdd_d vss_d / DCAP64LVT
XXFILLER_164_192 vdd_d vss_d / DCAP64LVT
XXFILLER_164_256 vdd_d vss_d / DCAP64LVT
XXFILLER_164_320 vdd_d vss_d / DCAP64LVT
XXFILLER_164_384 vdd_d vss_d / DCAP64LVT
XXFILLER_164_448 vdd_d vss_d / DCAP64LVT
XXFILLER_164_512 vdd_d vss_d / DCAP64LVT
XXFILLER_164_576 vdd_d vss_d / DCAP64LVT
XXFILLER_164_640 vdd_d vss_d / DCAP64LVT
XXFILLER_164_704 vdd_d vss_d / DCAP64LVT
XXFILLER_164_768 vdd_d vss_d / DCAP64LVT
XXFILLER_164_832 vdd_d vss_d / DCAP64LVT
XXFILLER_164_896 vdd_d vss_d / DCAP64LVT
XXFILLER_164_960 vdd_d vss_d / DCAP64LVT
XXFILLER_164_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_164_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_164_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_164_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_164_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_164_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_164_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_164_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_164_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_164_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_164_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_164_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_164_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_164_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_164_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_164_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_164_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_164_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_164_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_164_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_165_0 vdd_d vss_d / DCAP64LVT
XXFILLER_165_64 vdd_d vss_d / DCAP64LVT
XXFILLER_165_128 vdd_d vss_d / DCAP64LVT
XXFILLER_165_192 vdd_d vss_d / DCAP64LVT
XXFILLER_165_256 vdd_d vss_d / DCAP64LVT
XXFILLER_165_320 vdd_d vss_d / DCAP64LVT
XXFILLER_165_384 vdd_d vss_d / DCAP64LVT
XXFILLER_165_448 vdd_d vss_d / DCAP64LVT
XXFILLER_165_512 vdd_d vss_d / DCAP64LVT
XXFILLER_165_576 vdd_d vss_d / DCAP64LVT
XXFILLER_165_640 vdd_d vss_d / DCAP64LVT
XXFILLER_165_704 vdd_d vss_d / DCAP64LVT
XXFILLER_165_768 vdd_d vss_d / DCAP64LVT
XXFILLER_165_832 vdd_d vss_d / DCAP64LVT
XXFILLER_165_896 vdd_d vss_d / DCAP64LVT
XXFILLER_165_960 vdd_d vss_d / DCAP64LVT
XXFILLER_165_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_165_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_165_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_165_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_165_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_165_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_165_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_165_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_165_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_165_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_165_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_165_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_165_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_165_1889 vdd_d vss_d / DCAP64LVT
XXFILLER_165_1953 vdd_d vss_d / DCAP64LVT
XXFILLER_165_2017 vdd_d vss_d / DCAP64LVT
XXFILLER_165_2081 vdd_d vss_d / DCAP64LVT
XXFILLER_165_2145 vdd_d vss_d / DCAP64LVT
XXFILLER_165_2209 vdd_d vss_d / DCAP64LVT
XXFILLER_165_2273 vdd_d vss_d / DCAP64LVT
XXFILLER_166_0 vdd_d vss_d / DCAP64LVT
XXFILLER_166_64 vdd_d vss_d / DCAP64LVT
XXFILLER_166_128 vdd_d vss_d / DCAP64LVT
XXFILLER_166_192 vdd_d vss_d / DCAP64LVT
XXFILLER_166_256 vdd_d vss_d / DCAP64LVT
XXFILLER_166_320 vdd_d vss_d / DCAP64LVT
XXFILLER_166_384 vdd_d vss_d / DCAP64LVT
XXFILLER_166_448 vdd_d vss_d / DCAP64LVT
XXFILLER_166_512 vdd_d vss_d / DCAP64LVT
XXFILLER_166_576 vdd_d vss_d / DCAP64LVT
XXFILLER_166_640 vdd_d vss_d / DCAP64LVT
XXFILLER_166_704 vdd_d vss_d / DCAP64LVT
XXFILLER_166_768 vdd_d vss_d / DCAP64LVT
XXFILLER_166_832 vdd_d vss_d / DCAP64LVT
XXFILLER_166_942 vdd_d vss_d / DCAP64LVT
XXFILLER_166_1006 vdd_d vss_d / DCAP64LVT
XXFILLER_166_1070 vdd_d vss_d / DCAP64LVT
XXFILLER_166_1134 vdd_d vss_d / DCAP64LVT
XXFILLER_166_1198 vdd_d vss_d / DCAP64LVT
XXFILLER_166_1262 vdd_d vss_d / DCAP64LVT
XXFILLER_166_1326 vdd_d vss_d / DCAP64LVT
XXFILLER_166_1443 vdd_d vss_d / DCAP64LVT
XXFILLER_166_1507 vdd_d vss_d / DCAP64LVT
XXFILLER_166_1571 vdd_d vss_d / DCAP64LVT
XXFILLER_166_1635 vdd_d vss_d / DCAP64LVT
XXFILLER_166_1699 vdd_d vss_d / DCAP64LVT
XXFILLER_166_1763 vdd_d vss_d / DCAP64LVT
XXFILLER_166_1900 vdd_d vss_d / DCAP64LVT
XXFILLER_166_1964 vdd_d vss_d / DCAP64LVT
XXFILLER_166_2028 vdd_d vss_d / DCAP64LVT
XXFILLER_166_2092 vdd_d vss_d / DCAP64LVT
XXFILLER_166_2156 vdd_d vss_d / DCAP64LVT
XXFILLER_166_2220 vdd_d vss_d / DCAP64LVT
XXFILLER_166_2284 vdd_d vss_d / DCAP64LVT
XXFILLER_167_0 vdd_d vss_d / DCAP64LVT
XXFILLER_167_64 vdd_d vss_d / DCAP64LVT
XXFILLER_167_128 vdd_d vss_d / DCAP64LVT
XXFILLER_167_192 vdd_d vss_d / DCAP64LVT
XXFILLER_167_587 vdd_d vss_d / DCAP64LVT
XXFILLER_167_651 vdd_d vss_d / DCAP64LVT
XXFILLER_167_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_167_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_167_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_167_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_167_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_167_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_167_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_167_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_168_0 vdd_d vss_d / DCAP64LVT
XXFILLER_168_64 vdd_d vss_d / DCAP64LVT
XXFILLER_168_128 vdd_d vss_d / DCAP64LVT
XXFILLER_168_192 vdd_d vss_d / DCAP64LVT
XXFILLER_168_587 vdd_d vss_d / DCAP64LVT
XXFILLER_168_651 vdd_d vss_d / DCAP64LVT
XXFILLER_168_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_168_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_168_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_168_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_168_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_168_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_168_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_168_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_169_0 vdd_d vss_d / DCAP64LVT
XXFILLER_169_64 vdd_d vss_d / DCAP64LVT
XXFILLER_169_128 vdd_d vss_d / DCAP64LVT
XXFILLER_169_192 vdd_d vss_d / DCAP64LVT
XXFILLER_169_587 vdd_d vss_d / DCAP64LVT
XXFILLER_169_651 vdd_d vss_d / DCAP64LVT
XXFILLER_169_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_169_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_169_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_169_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_169_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_169_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_169_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_169_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_170_0 vdd_d vss_d / DCAP64LVT
XXFILLER_170_64 vdd_d vss_d / DCAP64LVT
XXFILLER_170_128 vdd_d vss_d / DCAP64LVT
XXFILLER_170_192 vdd_d vss_d / DCAP64LVT
XXFILLER_170_587 vdd_d vss_d / DCAP64LVT
XXFILLER_170_651 vdd_d vss_d / DCAP64LVT
XXFILLER_170_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_170_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_170_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_170_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_170_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_170_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_170_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_170_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_171_0 vdd_d vss_d / DCAP64LVT
XXFILLER_171_64 vdd_d vss_d / DCAP64LVT
XXFILLER_171_128 vdd_d vss_d / DCAP64LVT
XXFILLER_171_192 vdd_d vss_d / DCAP64LVT
XXFILLER_171_587 vdd_d vss_d / DCAP64LVT
XXFILLER_171_651 vdd_d vss_d / DCAP64LVT
XXFILLER_171_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_171_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_171_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_171_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_171_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_171_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_171_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_171_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_172_0 vdd_d vss_d / DCAP64LVT
XXFILLER_172_64 vdd_d vss_d / DCAP64LVT
XXFILLER_172_128 vdd_d vss_d / DCAP64LVT
XXFILLER_172_192 vdd_d vss_d / DCAP64LVT
XXFILLER_172_587 vdd_d vss_d / DCAP64LVT
XXFILLER_172_651 vdd_d vss_d / DCAP64LVT
XXFILLER_172_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_172_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_172_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_172_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_172_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_172_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_172_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_172_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_173_0 vdd_d vss_d / DCAP64LVT
XXFILLER_173_64 vdd_d vss_d / DCAP64LVT
XXFILLER_173_128 vdd_d vss_d / DCAP64LVT
XXFILLER_173_192 vdd_d vss_d / DCAP64LVT
XXFILLER_173_587 vdd_d vss_d / DCAP64LVT
XXFILLER_173_651 vdd_d vss_d / DCAP64LVT
XXFILLER_173_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_173_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_173_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_173_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_173_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_173_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_173_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_173_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_174_0 vdd_d vss_d / DCAP64LVT
XXFILLER_174_64 vdd_d vss_d / DCAP64LVT
XXFILLER_174_128 vdd_d vss_d / DCAP64LVT
XXFILLER_174_192 vdd_d vss_d / DCAP64LVT
XXFILLER_174_587 vdd_d vss_d / DCAP64LVT
XXFILLER_174_651 vdd_d vss_d / DCAP64LVT
XXFILLER_174_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_174_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_174_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_174_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_174_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_174_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_174_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_174_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_175_0 vdd_d vss_d / DCAP64LVT
XXFILLER_175_64 vdd_d vss_d / DCAP64LVT
XXFILLER_175_128 vdd_d vss_d / DCAP64LVT
XXFILLER_175_192 vdd_d vss_d / DCAP64LVT
XXFILLER_175_587 vdd_d vss_d / DCAP64LVT
XXFILLER_175_651 vdd_d vss_d / DCAP64LVT
XXFILLER_175_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_175_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_175_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_175_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_175_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_175_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_175_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_175_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_176_0 vdd_d vss_d / DCAP64LVT
XXFILLER_176_64 vdd_d vss_d / DCAP64LVT
XXFILLER_176_128 vdd_d vss_d / DCAP64LVT
XXFILLER_176_192 vdd_d vss_d / DCAP64LVT
XXFILLER_176_587 vdd_d vss_d / DCAP64LVT
XXFILLER_176_651 vdd_d vss_d / DCAP64LVT
XXFILLER_176_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_176_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_176_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_176_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_176_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_176_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_176_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_176_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_177_0 vdd_d vss_d / DCAP64LVT
XXFILLER_177_64 vdd_d vss_d / DCAP64LVT
XXFILLER_177_128 vdd_d vss_d / DCAP64LVT
XXFILLER_177_192 vdd_d vss_d / DCAP64LVT
XXFILLER_177_587 vdd_d vss_d / DCAP64LVT
XXFILLER_177_651 vdd_d vss_d / DCAP64LVT
XXFILLER_177_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_177_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_177_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_177_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_177_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_177_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_177_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_177_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_178_0 vdd_d vss_d / DCAP64LVT
XXFILLER_178_64 vdd_d vss_d / DCAP64LVT
XXFILLER_178_128 vdd_d vss_d / DCAP64LVT
XXFILLER_178_192 vdd_d vss_d / DCAP64LVT
XXFILLER_178_587 vdd_d vss_d / DCAP64LVT
XXFILLER_178_651 vdd_d vss_d / DCAP64LVT
XXFILLER_178_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_178_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_178_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_178_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_178_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_178_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_178_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_178_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_179_0 vdd_d vss_d / DCAP64LVT
XXFILLER_179_64 vdd_d vss_d / DCAP64LVT
XXFILLER_179_128 vdd_d vss_d / DCAP64LVT
XXFILLER_179_192 vdd_d vss_d / DCAP64LVT
XXFILLER_179_587 vdd_d vss_d / DCAP64LVT
XXFILLER_179_651 vdd_d vss_d / DCAP64LVT
XXFILLER_179_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_179_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_179_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_179_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_179_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_179_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_179_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_179_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_180_0 vdd_d vss_d / DCAP64LVT
XXFILLER_180_64 vdd_d vss_d / DCAP64LVT
XXFILLER_180_128 vdd_d vss_d / DCAP64LVT
XXFILLER_180_192 vdd_d vss_d / DCAP64LVT
XXFILLER_180_587 vdd_d vss_d / DCAP64LVT
XXFILLER_180_651 vdd_d vss_d / DCAP64LVT
XXFILLER_180_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_180_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_180_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_180_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_180_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_180_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_180_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_181_0 vdd_d vss_d / DCAP64LVT
XXFILLER_181_64 vdd_d vss_d / DCAP64LVT
XXFILLER_181_128 vdd_d vss_d / DCAP64LVT
XXFILLER_181_192 vdd_d vss_d / DCAP64LVT
XXFILLER_181_587 vdd_d vss_d / DCAP64LVT
XXFILLER_181_651 vdd_d vss_d / DCAP64LVT
XXFILLER_181_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_181_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_181_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_181_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_181_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_181_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_182_0 vdd_d vss_d / DCAP64LVT
XXFILLER_182_64 vdd_d vss_d / DCAP64LVT
XXFILLER_182_128 vdd_d vss_d / DCAP64LVT
XXFILLER_182_192 vdd_d vss_d / DCAP64LVT
XXFILLER_182_587 vdd_d vss_d / DCAP64LVT
XXFILLER_182_651 vdd_d vss_d / DCAP64LVT
XXFILLER_182_1105 vdd_d vss_d / DCAP64LVT
XXFILLER_182_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_182_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_182_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_182_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_182_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_182_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_183_0 vdd_d vss_d / DCAP64LVT
XXFILLER_183_64 vdd_d vss_d / DCAP64LVT
XXFILLER_183_128 vdd_d vss_d / DCAP64LVT
XXFILLER_183_192 vdd_d vss_d / DCAP64LVT
XXFILLER_183_587 vdd_d vss_d / DCAP64LVT
XXFILLER_183_651 vdd_d vss_d / DCAP64LVT
XXFILLER_183_1096 vdd_d vss_d / DCAP64LVT
XXFILLER_183_1160 vdd_d vss_d / DCAP64LVT
XXFILLER_183_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_183_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_183_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_183_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_183_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_183_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_184_0 vdd_d vss_d / DCAP64LVT
XXFILLER_184_64 vdd_d vss_d / DCAP64LVT
XXFILLER_184_128 vdd_d vss_d / DCAP64LVT
XXFILLER_184_192 vdd_d vss_d / DCAP64LVT
XXFILLER_184_587 vdd_d vss_d / DCAP64LVT
XXFILLER_184_651 vdd_d vss_d / DCAP64LVT
XXFILLER_184_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_184_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_184_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_184_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_184_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_184_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_184_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_184_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_185_0 vdd_d vss_d / DCAP64LVT
XXFILLER_185_64 vdd_d vss_d / DCAP64LVT
XXFILLER_185_128 vdd_d vss_d / DCAP64LVT
XXFILLER_185_192 vdd_d vss_d / DCAP64LVT
XXFILLER_185_587 vdd_d vss_d / DCAP64LVT
XXFILLER_185_651 vdd_d vss_d / DCAP64LVT
XXFILLER_185_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_185_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_185_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_185_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_185_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_185_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_185_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_185_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_186_0 vdd_d vss_d / DCAP64LVT
XXFILLER_186_64 vdd_d vss_d / DCAP64LVT
XXFILLER_186_128 vdd_d vss_d / DCAP64LVT
XXFILLER_186_192 vdd_d vss_d / DCAP64LVT
XXFILLER_186_587 vdd_d vss_d / DCAP64LVT
XXFILLER_186_651 vdd_d vss_d / DCAP64LVT
XXFILLER_186_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_186_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_186_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_186_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_186_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_186_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_186_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_186_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_187_0 vdd_d vss_d / DCAP64LVT
XXFILLER_187_64 vdd_d vss_d / DCAP64LVT
XXFILLER_187_128 vdd_d vss_d / DCAP64LVT
XXFILLER_187_192 vdd_d vss_d / DCAP64LVT
XXFILLER_187_587 vdd_d vss_d / DCAP64LVT
XXFILLER_187_651 vdd_d vss_d / DCAP64LVT
XXFILLER_187_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_187_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_187_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_187_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_187_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_187_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_187_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_187_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_188_0 vdd_d vss_d / DCAP64LVT
XXFILLER_188_64 vdd_d vss_d / DCAP64LVT
XXFILLER_188_128 vdd_d vss_d / DCAP64LVT
XXFILLER_188_192 vdd_d vss_d / DCAP64LVT
XXFILLER_188_587 vdd_d vss_d / DCAP64LVT
XXFILLER_188_651 vdd_d vss_d / DCAP64LVT
XXFILLER_188_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_188_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_188_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_188_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_188_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_188_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_188_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_188_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_189_0 vdd_d vss_d / DCAP64LVT
XXFILLER_189_64 vdd_d vss_d / DCAP64LVT
XXFILLER_189_128 vdd_d vss_d / DCAP64LVT
XXFILLER_189_192 vdd_d vss_d / DCAP64LVT
XXFILLER_189_587 vdd_d vss_d / DCAP64LVT
XXFILLER_189_651 vdd_d vss_d / DCAP64LVT
XXFILLER_189_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_189_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_189_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_189_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_189_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_189_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_189_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_189_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_190_0 vdd_d vss_d / DCAP64LVT
XXFILLER_190_64 vdd_d vss_d / DCAP64LVT
XXFILLER_190_128 vdd_d vss_d / DCAP64LVT
XXFILLER_190_192 vdd_d vss_d / DCAP64LVT
XXFILLER_190_587 vdd_d vss_d / DCAP64LVT
XXFILLER_190_651 vdd_d vss_d / DCAP64LVT
XXFILLER_190_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_190_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_190_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_190_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_190_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_190_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_190_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_190_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_191_0 vdd_d vss_d / DCAP64LVT
XXFILLER_191_64 vdd_d vss_d / DCAP64LVT
XXFILLER_191_128 vdd_d vss_d / DCAP64LVT
XXFILLER_191_192 vdd_d vss_d / DCAP64LVT
XXFILLER_191_587 vdd_d vss_d / DCAP64LVT
XXFILLER_191_651 vdd_d vss_d / DCAP64LVT
XXFILLER_191_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_191_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_191_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_191_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_191_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_191_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_191_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_191_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_192_0 vdd_d vss_d / DCAP64LVT
XXFILLER_192_64 vdd_d vss_d / DCAP64LVT
XXFILLER_192_128 vdd_d vss_d / DCAP64LVT
XXFILLER_192_192 vdd_d vss_d / DCAP64LVT
XXFILLER_192_587 vdd_d vss_d / DCAP64LVT
XXFILLER_192_651 vdd_d vss_d / DCAP64LVT
XXFILLER_192_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_192_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_192_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_192_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_192_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_192_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_192_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_192_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_193_0 vdd_d vss_d / DCAP64LVT
XXFILLER_193_64 vdd_d vss_d / DCAP64LVT
XXFILLER_193_128 vdd_d vss_d / DCAP64LVT
XXFILLER_193_192 vdd_d vss_d / DCAP64LVT
XXFILLER_193_587 vdd_d vss_d / DCAP64LVT
XXFILLER_193_651 vdd_d vss_d / DCAP64LVT
XXFILLER_193_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_193_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_193_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_193_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_193_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_193_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_193_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_193_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_194_0 vdd_d vss_d / DCAP64LVT
XXFILLER_194_64 vdd_d vss_d / DCAP64LVT
XXFILLER_194_128 vdd_d vss_d / DCAP64LVT
XXFILLER_194_192 vdd_d vss_d / DCAP64LVT
XXFILLER_194_587 vdd_d vss_d / DCAP64LVT
XXFILLER_194_651 vdd_d vss_d / DCAP64LVT
XXFILLER_194_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_194_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_194_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_194_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_194_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_194_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_194_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_194_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_195_0 vdd_d vss_d / DCAP64LVT
XXFILLER_195_64 vdd_d vss_d / DCAP64LVT
XXFILLER_195_128 vdd_d vss_d / DCAP64LVT
XXFILLER_195_192 vdd_d vss_d / DCAP64LVT
XXFILLER_195_587 vdd_d vss_d / DCAP64LVT
XXFILLER_195_651 vdd_d vss_d / DCAP64LVT
XXFILLER_195_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_195_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_195_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_195_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_195_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_195_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_195_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_195_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_196_0 vdd_d vss_d / DCAP64LVT
XXFILLER_196_64 vdd_d vss_d / DCAP64LVT
XXFILLER_196_128 vdd_d vss_d / DCAP64LVT
XXFILLER_196_192 vdd_d vss_d / DCAP64LVT
XXFILLER_196_587 vdd_d vss_d / DCAP64LVT
XXFILLER_196_651 vdd_d vss_d / DCAP64LVT
XXFILLER_196_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_196_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_196_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_196_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_196_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_196_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_196_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_196_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_197_0 vdd_d vss_d / DCAP64LVT
XXFILLER_197_64 vdd_d vss_d / DCAP64LVT
XXFILLER_197_128 vdd_d vss_d / DCAP64LVT
XXFILLER_197_192 vdd_d vss_d / DCAP64LVT
XXFILLER_197_587 vdd_d vss_d / DCAP64LVT
XXFILLER_197_651 vdd_d vss_d / DCAP64LVT
XXFILLER_197_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_197_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_197_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_197_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_197_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_197_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_197_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_197_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_198_0 vdd_d vss_d / DCAP64LVT
XXFILLER_198_64 vdd_d vss_d / DCAP64LVT
XXFILLER_198_128 vdd_d vss_d / DCAP64LVT
XXFILLER_198_192 vdd_d vss_d / DCAP64LVT
XXFILLER_198_587 vdd_d vss_d / DCAP64LVT
XXFILLER_198_651 vdd_d vss_d / DCAP64LVT
XXFILLER_198_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_198_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_198_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_198_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_198_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_198_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_198_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_198_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_199_0 vdd_d vss_d / DCAP64LVT
XXFILLER_199_64 vdd_d vss_d / DCAP64LVT
XXFILLER_199_128 vdd_d vss_d / DCAP64LVT
XXFILLER_199_192 vdd_d vss_d / DCAP64LVT
XXFILLER_199_587 vdd_d vss_d / DCAP64LVT
XXFILLER_199_651 vdd_d vss_d / DCAP64LVT
XXFILLER_199_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_199_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_199_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_199_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_199_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_199_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_199_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_199_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_200_0 vdd_d vss_d / DCAP64LVT
XXFILLER_200_64 vdd_d vss_d / DCAP64LVT
XXFILLER_200_128 vdd_d vss_d / DCAP64LVT
XXFILLER_200_192 vdd_d vss_d / DCAP64LVT
XXFILLER_200_587 vdd_d vss_d / DCAP64LVT
XXFILLER_200_651 vdd_d vss_d / DCAP64LVT
XXFILLER_200_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_200_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_200_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_200_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_200_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_200_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_200_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_200_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_201_0 vdd_d vss_d / DCAP64LVT
XXFILLER_201_64 vdd_d vss_d / DCAP64LVT
XXFILLER_201_128 vdd_d vss_d / DCAP64LVT
XXFILLER_201_192 vdd_d vss_d / DCAP64LVT
XXFILLER_201_587 vdd_d vss_d / DCAP64LVT
XXFILLER_201_651 vdd_d vss_d / DCAP64LVT
XXFILLER_201_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_201_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_201_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_201_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_201_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_201_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_201_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_201_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_202_0 vdd_d vss_d / DCAP64LVT
XXFILLER_202_64 vdd_d vss_d / DCAP64LVT
XXFILLER_202_128 vdd_d vss_d / DCAP64LVT
XXFILLER_202_192 vdd_d vss_d / DCAP64LVT
XXFILLER_202_587 vdd_d vss_d / DCAP64LVT
XXFILLER_202_651 vdd_d vss_d / DCAP64LVT
XXFILLER_202_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_202_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_202_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_202_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_202_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_202_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_202_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_202_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_203_0 vdd_d vss_d / DCAP64LVT
XXFILLER_203_64 vdd_d vss_d / DCAP64LVT
XXFILLER_203_128 vdd_d vss_d / DCAP64LVT
XXFILLER_203_192 vdd_d vss_d / DCAP64LVT
XXFILLER_203_587 vdd_d vss_d / DCAP64LVT
XXFILLER_203_651 vdd_d vss_d / DCAP64LVT
XXFILLER_203_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_203_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_203_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_203_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_203_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_203_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_203_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_203_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_204_0 vdd_d vss_d / DCAP64LVT
XXFILLER_204_64 vdd_d vss_d / DCAP64LVT
XXFILLER_204_128 vdd_d vss_d / DCAP64LVT
XXFILLER_204_192 vdd_d vss_d / DCAP64LVT
XXFILLER_204_587 vdd_d vss_d / DCAP64LVT
XXFILLER_204_651 vdd_d vss_d / DCAP64LVT
XXFILLER_204_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_204_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_204_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_204_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_204_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_204_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_204_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_204_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_205_0 vdd_d vss_d / DCAP64LVT
XXFILLER_205_64 vdd_d vss_d / DCAP64LVT
XXFILLER_205_128 vdd_d vss_d / DCAP64LVT
XXFILLER_205_192 vdd_d vss_d / DCAP64LVT
XXFILLER_205_587 vdd_d vss_d / DCAP64LVT
XXFILLER_205_651 vdd_d vss_d / DCAP64LVT
XXFILLER_205_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_205_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_205_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_205_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_205_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_205_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_205_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_205_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_206_0 vdd_d vss_d / DCAP64LVT
XXFILLER_206_64 vdd_d vss_d / DCAP64LVT
XXFILLER_206_128 vdd_d vss_d / DCAP64LVT
XXFILLER_206_192 vdd_d vss_d / DCAP64LVT
XXFILLER_206_256 vdd_d vss_d / DCAP64LVT
XXFILLER_206_320 vdd_d vss_d / DCAP64LVT
XXFILLER_206_447 vdd_d vss_d / DCAP64LVT
XXFILLER_206_511 vdd_d vss_d / DCAP64LVT
XXFILLER_206_575 vdd_d vss_d / DCAP64LVT
XXFILLER_206_639 vdd_d vss_d / DCAP64LVT
XXFILLER_206_703 vdd_d vss_d / DCAP64LVT
XXFILLER_206_767 vdd_d vss_d / DCAP64LVT
XXFILLER_206_831 vdd_d vss_d / DCAP64LVT
XXFILLER_206_956 vdd_d vss_d / DCAP64LVT
XXFILLER_206_1020 vdd_d vss_d / DCAP64LVT
XXFILLER_206_1084 vdd_d vss_d / DCAP64LVT
XXFILLER_206_1148 vdd_d vss_d / DCAP64LVT
XXFILLER_206_1212 vdd_d vss_d / DCAP64LVT
XXFILLER_206_1276 vdd_d vss_d / DCAP64LVT
XXFILLER_206_1340 vdd_d vss_d / DCAP64LVT
XXFILLER_206_1444 vdd_d vss_d / DCAP64LVT
XXFILLER_206_1508 vdd_d vss_d / DCAP64LVT
XXFILLER_206_1572 vdd_d vss_d / DCAP64LVT
XXFILLER_206_1636 vdd_d vss_d / DCAP64LVT
XXFILLER_206_1700 vdd_d vss_d / DCAP64LVT
XXFILLER_206_1764 vdd_d vss_d / DCAP64LVT
XXFILLER_206_1828 vdd_d vss_d / DCAP64LVT
XXFILLER_206_1892 vdd_d vss_d / DCAP64LVT
XXFILLER_206_1956 vdd_d vss_d / DCAP64LVT
XXFILLER_206_2020 vdd_d vss_d / DCAP64LVT
XXFILLER_206_2084 vdd_d vss_d / DCAP64LVT
XXFILLER_206_2148 vdd_d vss_d / DCAP64LVT
XXFILLER_206_2212 vdd_d vss_d / DCAP64LVT
XXFILLER_206_2276 vdd_d vss_d / DCAP64LVT
XXFILLER_207_0 vdd_d vss_d / DCAP64LVT
XXFILLER_207_64 vdd_d vss_d / DCAP64LVT
XXFILLER_207_128 vdd_d vss_d / DCAP64LVT
XXFILLER_207_192 vdd_d vss_d / DCAP64LVT
XXFILLER_207_256 vdd_d vss_d / DCAP64LVT
XXFILLER_207_320 vdd_d vss_d / DCAP64LVT
XXFILLER_207_384 vdd_d vss_d / DCAP64LVT
XXFILLER_207_448 vdd_d vss_d / DCAP64LVT
XXFILLER_207_512 vdd_d vss_d / DCAP64LVT
XXFILLER_207_576 vdd_d vss_d / DCAP64LVT
XXFILLER_207_640 vdd_d vss_d / DCAP64LVT
XXFILLER_207_704 vdd_d vss_d / DCAP64LVT
XXFILLER_207_768 vdd_d vss_d / DCAP64LVT
XXFILLER_207_832 vdd_d vss_d / DCAP64LVT
XXFILLER_207_950 vdd_d vss_d / DCAP64LVT
XXFILLER_207_1014 vdd_d vss_d / DCAP64LVT
XXFILLER_207_1078 vdd_d vss_d / DCAP64LVT
XXFILLER_207_1142 vdd_d vss_d / DCAP64LVT
XXFILLER_207_1206 vdd_d vss_d / DCAP64LVT
XXFILLER_207_1270 vdd_d vss_d / DCAP64LVT
XXFILLER_207_1334 vdd_d vss_d / DCAP64LVT
XXFILLER_207_1398 vdd_d vss_d / DCAP64LVT
XXFILLER_207_1462 vdd_d vss_d / DCAP64LVT
XXFILLER_207_1526 vdd_d vss_d / DCAP64LVT
XXFILLER_207_1590 vdd_d vss_d / DCAP64LVT
XXFILLER_207_1654 vdd_d vss_d / DCAP64LVT
XXFILLER_207_1718 vdd_d vss_d / DCAP64LVT
XXFILLER_207_1782 vdd_d vss_d / DCAP64LVT
XXFILLER_207_1846 vdd_d vss_d / DCAP64LVT
XXFILLER_207_1910 vdd_d vss_d / DCAP64LVT
XXFILLER_207_1974 vdd_d vss_d / DCAP64LVT
XXFILLER_207_2038 vdd_d vss_d / DCAP64LVT
XXFILLER_207_2102 vdd_d vss_d / DCAP64LVT
XXFILLER_207_2166 vdd_d vss_d / DCAP64LVT
XXFILLER_207_2230 vdd_d vss_d / DCAP64LVT
XXFILLER_208_0 vdd_d vss_d / DCAP64LVT
XXFILLER_208_64 vdd_d vss_d / DCAP64LVT
XXFILLER_208_128 vdd_d vss_d / DCAP64LVT
XXFILLER_208_192 vdd_d vss_d / DCAP64LVT
XXFILLER_208_256 vdd_d vss_d / DCAP64LVT
XXFILLER_208_320 vdd_d vss_d / DCAP64LVT
XXFILLER_208_384 vdd_d vss_d / DCAP64LVT
XXFILLER_208_448 vdd_d vss_d / DCAP64LVT
XXFILLER_208_512 vdd_d vss_d / DCAP64LVT
XXFILLER_208_576 vdd_d vss_d / DCAP64LVT
XXFILLER_208_640 vdd_d vss_d / DCAP64LVT
XXFILLER_208_704 vdd_d vss_d / DCAP64LVT
XXFILLER_208_768 vdd_d vss_d / DCAP64LVT
XXFILLER_208_832 vdd_d vss_d / DCAP64LVT
XXFILLER_208_896 vdd_d vss_d / DCAP64LVT
XXFILLER_208_960 vdd_d vss_d / DCAP64LVT
XXFILLER_208_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_208_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_208_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_208_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_208_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_208_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_208_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_208_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_208_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_208_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_208_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_208_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_208_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_208_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_208_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_208_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_208_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_208_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_208_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_208_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_209_0 vdd_d vss_d / DCAP64LVT
XXFILLER_209_64 vdd_d vss_d / DCAP64LVT
XXFILLER_209_128 vdd_d vss_d / DCAP64LVT
XXFILLER_209_192 vdd_d vss_d / DCAP64LVT
XXFILLER_209_256 vdd_d vss_d / DCAP64LVT
XXFILLER_209_320 vdd_d vss_d / DCAP64LVT
XXFILLER_209_384 vdd_d vss_d / DCAP64LVT
XXFILLER_209_448 vdd_d vss_d / DCAP64LVT
XXFILLER_209_512 vdd_d vss_d / DCAP64LVT
XXFILLER_209_576 vdd_d vss_d / DCAP64LVT
XXFILLER_209_640 vdd_d vss_d / DCAP64LVT
XXFILLER_209_704 vdd_d vss_d / DCAP64LVT
XXFILLER_209_768 vdd_d vss_d / DCAP64LVT
XXFILLER_209_832 vdd_d vss_d / DCAP64LVT
XXFILLER_209_896 vdd_d vss_d / DCAP64LVT
XXFILLER_209_960 vdd_d vss_d / DCAP64LVT
XXFILLER_209_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_209_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_209_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_209_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_209_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_209_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_209_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_209_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_209_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_209_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_209_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_209_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_209_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_209_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_209_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_209_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_209_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_209_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_209_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_209_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_210_0 vdd_d vss_d / DCAP64LVT
XXFILLER_210_64 vdd_d vss_d / DCAP64LVT
XXFILLER_210_128 vdd_d vss_d / DCAP64LVT
XXFILLER_210_192 vdd_d vss_d / DCAP64LVT
XXFILLER_210_256 vdd_d vss_d / DCAP64LVT
XXFILLER_210_320 vdd_d vss_d / DCAP64LVT
XXFILLER_210_384 vdd_d vss_d / DCAP64LVT
XXFILLER_210_448 vdd_d vss_d / DCAP64LVT
XXFILLER_210_512 vdd_d vss_d / DCAP64LVT
XXFILLER_210_576 vdd_d vss_d / DCAP64LVT
XXFILLER_210_640 vdd_d vss_d / DCAP64LVT
XXFILLER_210_704 vdd_d vss_d / DCAP64LVT
XXFILLER_210_768 vdd_d vss_d / DCAP64LVT
XXFILLER_210_832 vdd_d vss_d / DCAP64LVT
XXFILLER_210_896 vdd_d vss_d / DCAP64LVT
XXFILLER_210_960 vdd_d vss_d / DCAP64LVT
XXFILLER_210_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_210_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_210_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_210_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_210_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_210_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_210_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_210_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_210_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_210_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_210_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_210_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_210_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_210_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_210_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_210_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_210_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_210_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_210_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_210_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_211_0 vdd_d vss_d / DCAP64LVT
XXFILLER_211_64 vdd_d vss_d / DCAP64LVT
XXFILLER_211_128 vdd_d vss_d / DCAP64LVT
XXFILLER_211_192 vdd_d vss_d / DCAP64LVT
XXFILLER_211_256 vdd_d vss_d / DCAP64LVT
XXFILLER_211_320 vdd_d vss_d / DCAP64LVT
XXFILLER_211_384 vdd_d vss_d / DCAP64LVT
XXFILLER_211_448 vdd_d vss_d / DCAP64LVT
XXFILLER_211_512 vdd_d vss_d / DCAP64LVT
XXFILLER_211_576 vdd_d vss_d / DCAP64LVT
XXFILLER_211_640 vdd_d vss_d / DCAP64LVT
XXFILLER_211_704 vdd_d vss_d / DCAP64LVT
XXFILLER_211_768 vdd_d vss_d / DCAP64LVT
XXFILLER_211_832 vdd_d vss_d / DCAP64LVT
XXFILLER_211_896 vdd_d vss_d / DCAP64LVT
XXFILLER_211_960 vdd_d vss_d / DCAP64LVT
XXFILLER_211_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_211_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_211_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_211_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_211_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_211_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_211_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_211_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_211_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_211_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_211_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_211_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_211_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_211_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_211_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_211_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_211_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_211_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_211_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_211_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_212_0 vdd_d vss_d / DCAP64LVT
XXFILLER_212_64 vdd_d vss_d / DCAP64LVT
XXFILLER_212_128 vdd_d vss_d / DCAP64LVT
XXFILLER_212_192 vdd_d vss_d / DCAP64LVT
XXFILLER_212_256 vdd_d vss_d / DCAP64LVT
XXFILLER_212_320 vdd_d vss_d / DCAP64LVT
XXFILLER_212_384 vdd_d vss_d / DCAP64LVT
XXFILLER_212_448 vdd_d vss_d / DCAP64LVT
XXFILLER_212_512 vdd_d vss_d / DCAP64LVT
XXFILLER_212_576 vdd_d vss_d / DCAP64LVT
XXFILLER_212_640 vdd_d vss_d / DCAP64LVT
XXFILLER_212_704 vdd_d vss_d / DCAP64LVT
XXFILLER_212_768 vdd_d vss_d / DCAP64LVT
XXFILLER_212_832 vdd_d vss_d / DCAP64LVT
XXFILLER_212_896 vdd_d vss_d / DCAP64LVT
XXFILLER_212_960 vdd_d vss_d / DCAP64LVT
XXFILLER_212_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_212_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_212_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_212_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_212_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_212_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_212_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_212_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_212_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_212_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_212_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_212_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_212_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_212_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_212_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_212_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_212_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_212_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_212_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_212_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_213_0 vdd_d vss_d / DCAP64LVT
XXFILLER_213_64 vdd_d vss_d / DCAP64LVT
XXFILLER_213_128 vdd_d vss_d / DCAP64LVT
XXFILLER_213_192 vdd_d vss_d / DCAP64LVT
XXFILLER_213_256 vdd_d vss_d / DCAP64LVT
XXFILLER_213_320 vdd_d vss_d / DCAP64LVT
XXFILLER_213_384 vdd_d vss_d / DCAP64LVT
XXFILLER_213_448 vdd_d vss_d / DCAP64LVT
XXFILLER_213_512 vdd_d vss_d / DCAP64LVT
XXFILLER_213_576 vdd_d vss_d / DCAP64LVT
XXFILLER_213_640 vdd_d vss_d / DCAP64LVT
XXFILLER_213_704 vdd_d vss_d / DCAP64LVT
XXFILLER_213_768 vdd_d vss_d / DCAP64LVT
XXFILLER_213_832 vdd_d vss_d / DCAP64LVT
XXFILLER_213_896 vdd_d vss_d / DCAP64LVT
XXFILLER_213_960 vdd_d vss_d / DCAP64LVT
XXFILLER_213_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_213_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_213_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_213_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_213_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_213_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_213_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_213_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_213_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_213_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_213_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_213_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_213_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_213_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_213_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_213_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_213_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_213_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_213_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_213_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_214_0 vdd_d vss_d / DCAP64LVT
XXFILLER_214_64 vdd_d vss_d / DCAP64LVT
XXFILLER_214_128 vdd_d vss_d / DCAP64LVT
XXFILLER_214_192 vdd_d vss_d / DCAP64LVT
XXFILLER_214_256 vdd_d vss_d / DCAP64LVT
XXFILLER_214_320 vdd_d vss_d / DCAP64LVT
XXFILLER_214_384 vdd_d vss_d / DCAP64LVT
XXFILLER_214_448 vdd_d vss_d / DCAP64LVT
XXFILLER_214_512 vdd_d vss_d / DCAP64LVT
XXFILLER_214_576 vdd_d vss_d / DCAP64LVT
XXFILLER_214_709 vdd_d vss_d / DCAP64LVT
XXFILLER_214_773 vdd_d vss_d / DCAP64LVT
XXFILLER_214_837 vdd_d vss_d / DCAP64LVT
XXFILLER_214_901 vdd_d vss_d / DCAP64LVT
XXFILLER_214_965 vdd_d vss_d / DCAP64LVT
XXFILLER_214_1029 vdd_d vss_d / DCAP64LVT
XXFILLER_214_1093 vdd_d vss_d / DCAP64LVT
XXFILLER_214_1157 vdd_d vss_d / DCAP64LVT
XXFILLER_214_1221 vdd_d vss_d / DCAP64LVT
XXFILLER_214_1285 vdd_d vss_d / DCAP64LVT
XXFILLER_214_1349 vdd_d vss_d / DCAP64LVT
XXFILLER_214_1413 vdd_d vss_d / DCAP64LVT
XXFILLER_214_1477 vdd_d vss_d / DCAP64LVT
XXFILLER_214_1541 vdd_d vss_d / DCAP64LVT
XXFILLER_214_1605 vdd_d vss_d / DCAP64LVT
XXFILLER_214_1669 vdd_d vss_d / DCAP64LVT
XXFILLER_214_1733 vdd_d vss_d / DCAP64LVT
XXFILLER_214_1797 vdd_d vss_d / DCAP64LVT
XXFILLER_214_1861 vdd_d vss_d / DCAP64LVT
XXFILLER_214_1937 vdd_d vss_d / DCAP64LVT
XXFILLER_214_2001 vdd_d vss_d / DCAP64LVT
XXFILLER_214_2065 vdd_d vss_d / DCAP64LVT
XXFILLER_214_2129 vdd_d vss_d / DCAP64LVT
XXFILLER_214_2193 vdd_d vss_d / DCAP64LVT
XXFILLER_214_2257 vdd_d vss_d / DCAP64LVT
XXFILLER_215_0 vdd_d vss_d / DCAP64LVT
XXFILLER_215_64 vdd_d vss_d / DCAP64LVT
XXFILLER_215_128 vdd_d vss_d / DCAP64LVT
XXFILLER_215_192 vdd_d vss_d / DCAP64LVT
XXFILLER_215_256 vdd_d vss_d / DCAP64LVT
XXFILLER_215_320 vdd_d vss_d / DCAP64LVT
XXFILLER_215_384 vdd_d vss_d / DCAP64LVT
XXFILLER_215_448 vdd_d vss_d / DCAP64LVT
XXFILLER_215_512 vdd_d vss_d / DCAP64LVT
XXFILLER_215_576 vdd_d vss_d / DCAP64LVT
XXFILLER_215_640 vdd_d vss_d / DCAP64LVT
XXFILLER_215_704 vdd_d vss_d / DCAP64LVT
XXFILLER_215_768 vdd_d vss_d / DCAP64LVT
XXFILLER_215_832 vdd_d vss_d / DCAP64LVT
XXFILLER_215_896 vdd_d vss_d / DCAP64LVT
XXFILLER_215_960 vdd_d vss_d / DCAP64LVT
XXFILLER_215_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_215_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_215_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_215_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_215_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_215_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_215_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_215_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_215_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_215_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_215_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_215_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_215_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_215_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_215_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_215_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_215_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_215_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_215_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_215_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_216_0 vdd_d vss_d / DCAP64LVT
XXFILLER_216_64 vdd_d vss_d / DCAP64LVT
XXFILLER_216_128 vdd_d vss_d / DCAP64LVT
XXFILLER_216_192 vdd_d vss_d / DCAP64LVT
XXFILLER_216_256 vdd_d vss_d / DCAP64LVT
XXFILLER_216_320 vdd_d vss_d / DCAP64LVT
XXFILLER_216_384 vdd_d vss_d / DCAP64LVT
XXFILLER_216_448 vdd_d vss_d / DCAP64LVT
XXFILLER_216_512 vdd_d vss_d / DCAP64LVT
XXFILLER_216_576 vdd_d vss_d / DCAP64LVT
XXFILLER_216_640 vdd_d vss_d / DCAP64LVT
XXFILLER_216_704 vdd_d vss_d / DCAP64LVT
XXFILLER_216_768 vdd_d vss_d / DCAP64LVT
XXFILLER_216_832 vdd_d vss_d / DCAP64LVT
XXFILLER_216_896 vdd_d vss_d / DCAP64LVT
XXFILLER_216_960 vdd_d vss_d / DCAP64LVT
XXFILLER_216_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_216_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_216_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_216_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_216_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_216_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_216_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_216_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_216_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_216_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_216_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_216_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_216_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_216_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_216_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_216_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_216_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_216_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_216_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_216_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_217_0 vdd_d vss_d / DCAP64LVT
XXFILLER_217_64 vdd_d vss_d / DCAP64LVT
XXFILLER_217_128 vdd_d vss_d / DCAP64LVT
XXFILLER_217_192 vdd_d vss_d / DCAP64LVT
XXFILLER_217_256 vdd_d vss_d / DCAP64LVT
XXFILLER_217_320 vdd_d vss_d / DCAP64LVT
XXFILLER_217_384 vdd_d vss_d / DCAP64LVT
XXFILLER_217_448 vdd_d vss_d / DCAP64LVT
XXFILLER_217_512 vdd_d vss_d / DCAP64LVT
XXFILLER_217_576 vdd_d vss_d / DCAP64LVT
XXFILLER_217_640 vdd_d vss_d / DCAP64LVT
XXFILLER_217_704 vdd_d vss_d / DCAP64LVT
XXFILLER_217_768 vdd_d vss_d / DCAP64LVT
XXFILLER_217_832 vdd_d vss_d / DCAP64LVT
XXFILLER_217_896 vdd_d vss_d / DCAP64LVT
XXFILLER_217_960 vdd_d vss_d / DCAP64LVT
XXFILLER_217_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_217_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_217_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_217_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_217_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_217_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_217_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_217_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_217_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_217_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_217_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_217_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_217_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_217_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_217_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_217_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_217_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_217_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_217_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_217_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_218_0 vdd_d vss_d / DCAP64LVT
XXFILLER_218_64 vdd_d vss_d / DCAP64LVT
XXFILLER_218_128 vdd_d vss_d / DCAP64LVT
XXFILLER_218_192 vdd_d vss_d / DCAP64LVT
XXFILLER_218_256 vdd_d vss_d / DCAP64LVT
XXFILLER_218_320 vdd_d vss_d / DCAP64LVT
XXFILLER_218_384 vdd_d vss_d / DCAP64LVT
XXFILLER_218_448 vdd_d vss_d / DCAP64LVT
XXFILLER_218_512 vdd_d vss_d / DCAP64LVT
XXFILLER_218_576 vdd_d vss_d / DCAP64LVT
XXFILLER_218_640 vdd_d vss_d / DCAP64LVT
XXFILLER_218_704 vdd_d vss_d / DCAP64LVT
XXFILLER_218_768 vdd_d vss_d / DCAP64LVT
XXFILLER_218_832 vdd_d vss_d / DCAP64LVT
XXFILLER_218_896 vdd_d vss_d / DCAP64LVT
XXFILLER_218_960 vdd_d vss_d / DCAP64LVT
XXFILLER_218_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_218_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_218_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_218_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_218_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_218_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_218_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_218_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_218_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_218_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_218_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_218_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_218_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_218_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_218_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_218_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_218_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_218_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_218_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_218_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_219_0 vdd_d vss_d / DCAP64LVT
XXFILLER_219_64 vdd_d vss_d / DCAP64LVT
XXFILLER_219_128 vdd_d vss_d / DCAP64LVT
XXFILLER_219_192 vdd_d vss_d / DCAP64LVT
XXFILLER_219_256 vdd_d vss_d / DCAP64LVT
XXFILLER_219_320 vdd_d vss_d / DCAP64LVT
XXFILLER_219_384 vdd_d vss_d / DCAP64LVT
XXFILLER_219_448 vdd_d vss_d / DCAP64LVT
XXFILLER_219_512 vdd_d vss_d / DCAP64LVT
XXFILLER_219_576 vdd_d vss_d / DCAP64LVT
XXFILLER_219_640 vdd_d vss_d / DCAP64LVT
XXFILLER_219_704 vdd_d vss_d / DCAP64LVT
XXFILLER_219_768 vdd_d vss_d / DCAP64LVT
XXFILLER_219_832 vdd_d vss_d / DCAP64LVT
XXFILLER_219_944 vdd_d vss_d / DCAP64LVT
XXFILLER_219_1008 vdd_d vss_d / DCAP64LVT
XXFILLER_219_1072 vdd_d vss_d / DCAP64LVT
XXFILLER_219_1136 vdd_d vss_d / DCAP64LVT
XXFILLER_219_1200 vdd_d vss_d / DCAP64LVT
XXFILLER_219_1264 vdd_d vss_d / DCAP64LVT
XXFILLER_219_1328 vdd_d vss_d / DCAP64LVT
XXFILLER_219_1392 vdd_d vss_d / DCAP64LVT
XXFILLER_219_1456 vdd_d vss_d / DCAP64LVT
XXFILLER_219_1520 vdd_d vss_d / DCAP64LVT
XXFILLER_219_1584 vdd_d vss_d / DCAP64LVT
XXFILLER_219_1648 vdd_d vss_d / DCAP64LVT
XXFILLER_219_1712 vdd_d vss_d / DCAP64LVT
XXFILLER_219_1776 vdd_d vss_d / DCAP64LVT
XXFILLER_219_1840 vdd_d vss_d / DCAP64LVT
XXFILLER_219_1904 vdd_d vss_d / DCAP64LVT
XXFILLER_219_1968 vdd_d vss_d / DCAP64LVT
XXFILLER_219_2032 vdd_d vss_d / DCAP64LVT
XXFILLER_219_2096 vdd_d vss_d / DCAP64LVT
XXFILLER_219_2160 vdd_d vss_d / DCAP64LVT
XXFILLER_219_2224 vdd_d vss_d / DCAP64LVT
XXFILLER_220_0 vdd_d vss_d / DCAP64LVT
XXFILLER_220_64 vdd_d vss_d / DCAP64LVT
XXFILLER_220_128 vdd_d vss_d / DCAP64LVT
XXFILLER_220_192 vdd_d vss_d / DCAP64LVT
XXFILLER_220_256 vdd_d vss_d / DCAP64LVT
XXFILLER_220_320 vdd_d vss_d / DCAP64LVT
XXFILLER_220_384 vdd_d vss_d / DCAP64LVT
XXFILLER_220_448 vdd_d vss_d / DCAP64LVT
XXFILLER_220_512 vdd_d vss_d / DCAP64LVT
XXFILLER_220_576 vdd_d vss_d / DCAP64LVT
XXFILLER_220_640 vdd_d vss_d / DCAP64LVT
XXFILLER_220_704 vdd_d vss_d / DCAP64LVT
XXFILLER_220_768 vdd_d vss_d / DCAP64LVT
XXFILLER_220_832 vdd_d vss_d / DCAP64LVT
XXFILLER_220_896 vdd_d vss_d / DCAP64LVT
XXFILLER_220_960 vdd_d vss_d / DCAP64LVT
XXFILLER_220_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_220_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_220_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_220_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_220_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_220_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_220_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_220_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_220_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_220_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_220_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_220_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_220_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_220_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_220_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_220_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_220_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_220_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_220_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_220_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_221_0 vdd_d vss_d / DCAP64LVT
XXFILLER_221_64 vdd_d vss_d / DCAP64LVT
XXFILLER_221_128 vdd_d vss_d / DCAP64LVT
XXFILLER_221_192 vdd_d vss_d / DCAP64LVT
XXFILLER_221_256 vdd_d vss_d / DCAP64LVT
XXFILLER_221_320 vdd_d vss_d / DCAP64LVT
XXFILLER_221_384 vdd_d vss_d / DCAP64LVT
XXFILLER_221_448 vdd_d vss_d / DCAP64LVT
XXFILLER_221_512 vdd_d vss_d / DCAP64LVT
XXFILLER_221_576 vdd_d vss_d / DCAP64LVT
XXFILLER_221_640 vdd_d vss_d / DCAP64LVT
XXFILLER_221_704 vdd_d vss_d / DCAP64LVT
XXFILLER_221_768 vdd_d vss_d / DCAP64LVT
XXFILLER_221_832 vdd_d vss_d / DCAP64LVT
XXFILLER_221_896 vdd_d vss_d / DCAP64LVT
XXFILLER_221_960 vdd_d vss_d / DCAP64LVT
XXFILLER_221_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_221_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_221_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_221_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_221_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_221_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_221_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_221_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_221_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_221_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_221_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_221_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_221_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_221_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_221_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_221_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_221_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_221_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_221_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_221_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_222_0 vdd_d vss_d / DCAP64LVT
XXFILLER_222_64 vdd_d vss_d / DCAP64LVT
XXFILLER_222_128 vdd_d vss_d / DCAP64LVT
XXFILLER_222_192 vdd_d vss_d / DCAP64LVT
XXFILLER_222_256 vdd_d vss_d / DCAP64LVT
XXFILLER_222_320 vdd_d vss_d / DCAP64LVT
XXFILLER_222_384 vdd_d vss_d / DCAP64LVT
XXFILLER_222_448 vdd_d vss_d / DCAP64LVT
XXFILLER_222_512 vdd_d vss_d / DCAP64LVT
XXFILLER_222_576 vdd_d vss_d / DCAP64LVT
XXFILLER_222_640 vdd_d vss_d / DCAP64LVT
XXFILLER_222_704 vdd_d vss_d / DCAP64LVT
XXFILLER_222_768 vdd_d vss_d / DCAP64LVT
XXFILLER_222_832 vdd_d vss_d / DCAP64LVT
XXFILLER_222_896 vdd_d vss_d / DCAP64LVT
XXFILLER_222_960 vdd_d vss_d / DCAP64LVT
XXFILLER_222_1024 vdd_d vss_d / DCAP64LVT
XXFILLER_222_1088 vdd_d vss_d / DCAP64LVT
XXFILLER_222_1152 vdd_d vss_d / DCAP64LVT
XXFILLER_222_1216 vdd_d vss_d / DCAP64LVT
XXFILLER_222_1280 vdd_d vss_d / DCAP64LVT
XXFILLER_222_1344 vdd_d vss_d / DCAP64LVT
XXFILLER_222_1408 vdd_d vss_d / DCAP64LVT
XXFILLER_222_1472 vdd_d vss_d / DCAP64LVT
XXFILLER_222_1536 vdd_d vss_d / DCAP64LVT
XXFILLER_222_1600 vdd_d vss_d / DCAP64LVT
XXFILLER_222_1664 vdd_d vss_d / DCAP64LVT
XXFILLER_222_1728 vdd_d vss_d / DCAP64LVT
XXFILLER_222_1792 vdd_d vss_d / DCAP64LVT
XXFILLER_222_1856 vdd_d vss_d / DCAP64LVT
XXFILLER_222_1920 vdd_d vss_d / DCAP64LVT
XXFILLER_222_1984 vdd_d vss_d / DCAP64LVT
XXFILLER_222_2048 vdd_d vss_d / DCAP64LVT
XXFILLER_222_2112 vdd_d vss_d / DCAP64LVT
XXFILLER_222_2176 vdd_d vss_d / DCAP64LVT
XXFILLER_222_2240 vdd_d vss_d / DCAP64LVT
XXFILLER_223_0 vdd_d vss_d / DCAP64LVT
XXFILLER_223_64 vdd_d vss_d / DCAP64LVT
XXFILLER_223_128 vdd_d vss_d / DCAP64LVT
XXFILLER_223_192 vdd_d vss_d / DCAP64LVT
XXFILLER_223_587 vdd_d vss_d / DCAP64LVT
XXFILLER_223_651 vdd_d vss_d / DCAP64LVT
XXFILLER_223_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_223_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_223_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_223_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_223_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_223_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_223_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_223_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_224_0 vdd_d vss_d / DCAP64LVT
XXFILLER_224_64 vdd_d vss_d / DCAP64LVT
XXFILLER_224_128 vdd_d vss_d / DCAP64LVT
XXFILLER_224_192 vdd_d vss_d / DCAP64LVT
XXFILLER_224_587 vdd_d vss_d / DCAP64LVT
XXFILLER_224_651 vdd_d vss_d / DCAP64LVT
XXFILLER_224_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_224_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_224_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_224_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_224_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_224_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_224_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_224_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_225_0 vdd_d vss_d / DCAP64LVT
XXFILLER_225_64 vdd_d vss_d / DCAP64LVT
XXFILLER_225_128 vdd_d vss_d / DCAP64LVT
XXFILLER_225_192 vdd_d vss_d / DCAP64LVT
XXFILLER_225_587 vdd_d vss_d / DCAP64LVT
XXFILLER_225_651 vdd_d vss_d / DCAP64LVT
XXFILLER_225_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_225_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_225_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_225_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_225_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_225_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_225_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_225_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_226_0 vdd_d vss_d / DCAP64LVT
XXFILLER_226_64 vdd_d vss_d / DCAP64LVT
XXFILLER_226_128 vdd_d vss_d / DCAP64LVT
XXFILLER_226_192 vdd_d vss_d / DCAP64LVT
XXFILLER_226_587 vdd_d vss_d / DCAP64LVT
XXFILLER_226_651 vdd_d vss_d / DCAP64LVT
XXFILLER_226_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_226_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_226_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_226_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_226_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_226_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_226_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_226_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_227_0 vdd_d vss_d / DCAP64LVT
XXFILLER_227_64 vdd_d vss_d / DCAP64LVT
XXFILLER_227_128 vdd_d vss_d / DCAP64LVT
XXFILLER_227_192 vdd_d vss_d / DCAP64LVT
XXFILLER_227_587 vdd_d vss_d / DCAP64LVT
XXFILLER_227_651 vdd_d vss_d / DCAP64LVT
XXFILLER_227_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_227_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_227_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_227_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_227_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_227_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_227_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_227_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_228_0 vdd_d vss_d / DCAP64LVT
XXFILLER_228_64 vdd_d vss_d / DCAP64LVT
XXFILLER_228_128 vdd_d vss_d / DCAP64LVT
XXFILLER_228_192 vdd_d vss_d / DCAP64LVT
XXFILLER_228_587 vdd_d vss_d / DCAP64LVT
XXFILLER_228_651 vdd_d vss_d / DCAP64LVT
XXFILLER_228_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_228_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_228_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_228_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_228_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_228_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_228_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_228_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_229_0 vdd_d vss_d / DCAP64LVT
XXFILLER_229_64 vdd_d vss_d / DCAP64LVT
XXFILLER_229_128 vdd_d vss_d / DCAP64LVT
XXFILLER_229_192 vdd_d vss_d / DCAP64LVT
XXFILLER_229_587 vdd_d vss_d / DCAP64LVT
XXFILLER_229_651 vdd_d vss_d / DCAP64LVT
XXFILLER_229_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_229_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_229_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_229_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_229_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_229_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_229_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_229_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_230_0 vdd_d vss_d / DCAP64LVT
XXFILLER_230_64 vdd_d vss_d / DCAP64LVT
XXFILLER_230_128 vdd_d vss_d / DCAP64LVT
XXFILLER_230_192 vdd_d vss_d / DCAP64LVT
XXFILLER_230_587 vdd_d vss_d / DCAP64LVT
XXFILLER_230_651 vdd_d vss_d / DCAP64LVT
XXFILLER_230_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_230_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_230_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_230_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_230_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_230_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_230_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_230_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_231_0 vdd_d vss_d / DCAP64LVT
XXFILLER_231_64 vdd_d vss_d / DCAP64LVT
XXFILLER_231_128 vdd_d vss_d / DCAP64LVT
XXFILLER_231_192 vdd_d vss_d / DCAP64LVT
XXFILLER_231_587 vdd_d vss_d / DCAP64LVT
XXFILLER_231_651 vdd_d vss_d / DCAP64LVT
XXFILLER_231_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_231_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_231_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_231_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_231_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_231_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_231_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_231_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_232_0 vdd_d vss_d / DCAP64LVT
XXFILLER_232_64 vdd_d vss_d / DCAP64LVT
XXFILLER_232_128 vdd_d vss_d / DCAP64LVT
XXFILLER_232_192 vdd_d vss_d / DCAP64LVT
XXFILLER_232_587 vdd_d vss_d / DCAP64LVT
XXFILLER_232_651 vdd_d vss_d / DCAP64LVT
XXFILLER_232_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_232_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_232_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_232_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_232_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_232_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_232_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_232_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_233_0 vdd_d vss_d / DCAP64LVT
XXFILLER_233_64 vdd_d vss_d / DCAP64LVT
XXFILLER_233_128 vdd_d vss_d / DCAP64LVT
XXFILLER_233_192 vdd_d vss_d / DCAP64LVT
XXFILLER_233_587 vdd_d vss_d / DCAP64LVT
XXFILLER_233_651 vdd_d vss_d / DCAP64LVT
XXFILLER_233_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_233_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_233_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_233_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_233_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_233_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_233_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_233_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_234_0 vdd_d vss_d / DCAP64LVT
XXFILLER_234_64 vdd_d vss_d / DCAP64LVT
XXFILLER_234_128 vdd_d vss_d / DCAP64LVT
XXFILLER_234_192 vdd_d vss_d / DCAP64LVT
XXFILLER_234_587 vdd_d vss_d / DCAP64LVT
XXFILLER_234_651 vdd_d vss_d / DCAP64LVT
XXFILLER_234_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_234_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_234_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_234_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_234_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_234_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_234_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_234_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_235_0 vdd_d vss_d / DCAP64LVT
XXFILLER_235_64 vdd_d vss_d / DCAP64LVT
XXFILLER_235_128 vdd_d vss_d / DCAP64LVT
XXFILLER_235_192 vdd_d vss_d / DCAP64LVT
XXFILLER_235_587 vdd_d vss_d / DCAP64LVT
XXFILLER_235_651 vdd_d vss_d / DCAP64LVT
XXFILLER_235_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_235_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_235_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_235_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_235_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_235_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_235_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_235_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_236_0 vdd_d vss_d / DCAP64LVT
XXFILLER_236_64 vdd_d vss_d / DCAP64LVT
XXFILLER_236_128 vdd_d vss_d / DCAP64LVT
XXFILLER_236_192 vdd_d vss_d / DCAP64LVT
XXFILLER_236_587 vdd_d vss_d / DCAP64LVT
XXFILLER_236_651 vdd_d vss_d / DCAP64LVT
XXFILLER_236_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_236_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_236_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_236_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_236_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_236_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_236_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_236_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_237_0 vdd_d vss_d / DCAP64LVT
XXFILLER_237_64 vdd_d vss_d / DCAP64LVT
XXFILLER_237_128 vdd_d vss_d / DCAP64LVT
XXFILLER_237_192 vdd_d vss_d / DCAP64LVT
XXFILLER_237_587 vdd_d vss_d / DCAP64LVT
XXFILLER_237_651 vdd_d vss_d / DCAP64LVT
XXFILLER_237_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_237_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_237_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_237_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_237_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_237_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_237_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_237_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_238_0 vdd_d vss_d / DCAP64LVT
XXFILLER_238_64 vdd_d vss_d / DCAP64LVT
XXFILLER_238_128 vdd_d vss_d / DCAP64LVT
XXFILLER_238_192 vdd_d vss_d / DCAP64LVT
XXFILLER_238_587 vdd_d vss_d / DCAP64LVT
XXFILLER_238_651 vdd_d vss_d / DCAP64LVT
XXFILLER_238_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_238_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_238_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_238_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_238_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_238_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_238_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_238_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_239_0 vdd_d vss_d / DCAP64LVT
XXFILLER_239_64 vdd_d vss_d / DCAP64LVT
XXFILLER_239_128 vdd_d vss_d / DCAP64LVT
XXFILLER_239_192 vdd_d vss_d / DCAP64LVT
XXFILLER_239_587 vdd_d vss_d / DCAP64LVT
XXFILLER_239_651 vdd_d vss_d / DCAP64LVT
XXFILLER_239_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_239_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_239_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_239_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_239_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_239_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_239_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_239_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_240_0 vdd_d vss_d / DCAP64LVT
XXFILLER_240_64 vdd_d vss_d / DCAP64LVT
XXFILLER_240_128 vdd_d vss_d / DCAP64LVT
XXFILLER_240_192 vdd_d vss_d / DCAP64LVT
XXFILLER_240_587 vdd_d vss_d / DCAP64LVT
XXFILLER_240_651 vdd_d vss_d / DCAP64LVT
XXFILLER_240_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_240_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_240_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_240_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_240_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_240_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_240_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_240_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_241_0 vdd_d vss_d / DCAP64LVT
XXFILLER_241_64 vdd_d vss_d / DCAP64LVT
XXFILLER_241_128 vdd_d vss_d / DCAP64LVT
XXFILLER_241_192 vdd_d vss_d / DCAP64LVT
XXFILLER_241_587 vdd_d vss_d / DCAP64LVT
XXFILLER_241_651 vdd_d vss_d / DCAP64LVT
XXFILLER_241_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_241_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_241_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_241_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_241_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_241_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_241_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_241_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_242_0 vdd_d vss_d / DCAP64LVT
XXFILLER_242_64 vdd_d vss_d / DCAP64LVT
XXFILLER_242_128 vdd_d vss_d / DCAP64LVT
XXFILLER_242_192 vdd_d vss_d / DCAP64LVT
XXFILLER_242_587 vdd_d vss_d / DCAP64LVT
XXFILLER_242_651 vdd_d vss_d / DCAP64LVT
XXFILLER_242_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_242_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_242_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_242_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_242_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_242_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_242_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_242_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_243_0 vdd_d vss_d / DCAP64LVT
XXFILLER_243_64 vdd_d vss_d / DCAP64LVT
XXFILLER_243_128 vdd_d vss_d / DCAP64LVT
XXFILLER_243_192 vdd_d vss_d / DCAP64LVT
XXFILLER_243_587 vdd_d vss_d / DCAP64LVT
XXFILLER_243_651 vdd_d vss_d / DCAP64LVT
XXFILLER_243_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_243_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_243_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_243_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_243_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_243_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_243_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_243_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_244_0 vdd_d vss_d / DCAP64LVT
XXFILLER_244_64 vdd_d vss_d / DCAP64LVT
XXFILLER_244_128 vdd_d vss_d / DCAP64LVT
XXFILLER_244_192 vdd_d vss_d / DCAP64LVT
XXFILLER_244_587 vdd_d vss_d / DCAP64LVT
XXFILLER_244_651 vdd_d vss_d / DCAP64LVT
XXFILLER_244_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_244_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_244_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_244_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_244_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_244_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_244_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_244_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_245_0 vdd_d vss_d / DCAP64LVT
XXFILLER_245_64 vdd_d vss_d / DCAP64LVT
XXFILLER_245_128 vdd_d vss_d / DCAP64LVT
XXFILLER_245_192 vdd_d vss_d / DCAP64LVT
XXFILLER_245_587 vdd_d vss_d / DCAP64LVT
XXFILLER_245_651 vdd_d vss_d / DCAP64LVT
XXFILLER_245_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_245_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_245_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_245_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_245_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_245_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_245_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_245_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_246_0 vdd_d vss_d / DCAP64LVT
XXFILLER_246_64 vdd_d vss_d / DCAP64LVT
XXFILLER_246_128 vdd_d vss_d / DCAP64LVT
XXFILLER_246_192 vdd_d vss_d / DCAP64LVT
XXFILLER_246_587 vdd_d vss_d / DCAP64LVT
XXFILLER_246_651 vdd_d vss_d / DCAP64LVT
XXFILLER_246_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_246_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_246_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_246_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_246_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_246_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_246_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_246_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_247_0 vdd_d vss_d / DCAP64LVT
XXFILLER_247_64 vdd_d vss_d / DCAP64LVT
XXFILLER_247_128 vdd_d vss_d / DCAP64LVT
XXFILLER_247_192 vdd_d vss_d / DCAP64LVT
XXFILLER_247_587 vdd_d vss_d / DCAP64LVT
XXFILLER_247_651 vdd_d vss_d / DCAP64LVT
XXFILLER_247_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_247_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_247_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_247_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_247_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_247_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_247_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_247_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_248_0 vdd_d vss_d / DCAP64LVT
XXFILLER_248_64 vdd_d vss_d / DCAP64LVT
XXFILLER_248_128 vdd_d vss_d / DCAP64LVT
XXFILLER_248_192 vdd_d vss_d / DCAP64LVT
XXFILLER_248_587 vdd_d vss_d / DCAP64LVT
XXFILLER_248_651 vdd_d vss_d / DCAP64LVT
XXFILLER_248_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_248_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_248_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_248_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_248_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_248_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_248_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_248_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_249_0 vdd_d vss_d / DCAP64LVT
XXFILLER_249_64 vdd_d vss_d / DCAP64LVT
XXFILLER_249_128 vdd_d vss_d / DCAP64LVT
XXFILLER_249_192 vdd_d vss_d / DCAP64LVT
XXFILLER_249_587 vdd_d vss_d / DCAP64LVT
XXFILLER_249_651 vdd_d vss_d / DCAP64LVT
XXFILLER_249_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_249_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_249_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_249_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_249_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_249_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_249_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_249_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_250_0 vdd_d vss_d / DCAP64LVT
XXFILLER_250_64 vdd_d vss_d / DCAP64LVT
XXFILLER_250_128 vdd_d vss_d / DCAP64LVT
XXFILLER_250_192 vdd_d vss_d / DCAP64LVT
XXFILLER_250_587 vdd_d vss_d / DCAP64LVT
XXFILLER_250_651 vdd_d vss_d / DCAP64LVT
XXFILLER_250_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_250_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_250_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_250_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_250_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_250_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_250_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_250_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_251_0 vdd_d vss_d / DCAP64LVT
XXFILLER_251_64 vdd_d vss_d / DCAP64LVT
XXFILLER_251_128 vdd_d vss_d / DCAP64LVT
XXFILLER_251_192 vdd_d vss_d / DCAP64LVT
XXFILLER_251_587 vdd_d vss_d / DCAP64LVT
XXFILLER_251_651 vdd_d vss_d / DCAP64LVT
XXFILLER_251_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_251_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_251_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_251_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_251_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_251_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_251_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_251_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_252_0 vdd_d vss_d / DCAP64LVT
XXFILLER_252_64 vdd_d vss_d / DCAP64LVT
XXFILLER_252_128 vdd_d vss_d / DCAP64LVT
XXFILLER_252_192 vdd_d vss_d / DCAP64LVT
XXFILLER_252_587 vdd_d vss_d / DCAP64LVT
XXFILLER_252_651 vdd_d vss_d / DCAP64LVT
XXFILLER_252_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_252_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_252_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_252_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_252_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_252_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_252_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_252_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_253_0 vdd_d vss_d / DCAP64LVT
XXFILLER_253_64 vdd_d vss_d / DCAP64LVT
XXFILLER_253_128 vdd_d vss_d / DCAP64LVT
XXFILLER_253_192 vdd_d vss_d / DCAP64LVT
XXFILLER_253_587 vdd_d vss_d / DCAP64LVT
XXFILLER_253_651 vdd_d vss_d / DCAP64LVT
XXFILLER_253_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_253_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_253_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_253_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_253_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_253_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_253_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_253_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_254_0 vdd_d vss_d / DCAP64LVT
XXFILLER_254_64 vdd_d vss_d / DCAP64LVT
XXFILLER_254_128 vdd_d vss_d / DCAP64LVT
XXFILLER_254_192 vdd_d vss_d / DCAP64LVT
XXFILLER_254_587 vdd_d vss_d / DCAP64LVT
XXFILLER_254_651 vdd_d vss_d / DCAP64LVT
XXFILLER_254_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_254_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_254_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_254_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_254_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_254_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_254_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_254_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_255_0 vdd_d vss_d / DCAP64LVT
XXFILLER_255_64 vdd_d vss_d / DCAP64LVT
XXFILLER_255_128 vdd_d vss_d / DCAP64LVT
XXFILLER_255_192 vdd_d vss_d / DCAP64LVT
XXFILLER_255_587 vdd_d vss_d / DCAP64LVT
XXFILLER_255_651 vdd_d vss_d / DCAP64LVT
XXFILLER_255_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_255_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_255_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_255_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_255_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_255_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_255_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_255_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_256_0 vdd_d vss_d / DCAP64LVT
XXFILLER_256_64 vdd_d vss_d / DCAP64LVT
XXFILLER_256_128 vdd_d vss_d / DCAP64LVT
XXFILLER_256_192 vdd_d vss_d / DCAP64LVT
XXFILLER_256_587 vdd_d vss_d / DCAP64LVT
XXFILLER_256_651 vdd_d vss_d / DCAP64LVT
XXFILLER_256_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_256_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_256_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_256_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_256_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_256_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_256_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_256_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_257_0 vdd_d vss_d / DCAP64LVT
XXFILLER_257_64 vdd_d vss_d / DCAP64LVT
XXFILLER_257_128 vdd_d vss_d / DCAP64LVT
XXFILLER_257_192 vdd_d vss_d / DCAP64LVT
XXFILLER_257_587 vdd_d vss_d / DCAP64LVT
XXFILLER_257_651 vdd_d vss_d / DCAP64LVT
XXFILLER_257_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_257_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_257_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_257_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_257_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_257_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_257_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_257_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_258_0 vdd_d vss_d / DCAP64LVT
XXFILLER_258_64 vdd_d vss_d / DCAP64LVT
XXFILLER_258_128 vdd_d vss_d / DCAP64LVT
XXFILLER_258_192 vdd_d vss_d / DCAP64LVT
XXFILLER_258_587 vdd_d vss_d / DCAP64LVT
XXFILLER_258_651 vdd_d vss_d / DCAP64LVT
XXFILLER_258_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_258_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_258_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_258_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_258_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_258_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_258_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_258_2279 vdd_d vss_d / DCAP64LVT
XXFILLER_259_0 vdd_d vss_d / DCAP64LVT
XXFILLER_259_64 vdd_d vss_d / DCAP64LVT
XXFILLER_259_128 vdd_d vss_d / DCAP64LVT
XXFILLER_259_192 vdd_d vss_d / DCAP64LVT
XXFILLER_259_587 vdd_d vss_d / DCAP64LVT
XXFILLER_259_651 vdd_d vss_d / DCAP64LVT
XXFILLER_259_1087 vdd_d vss_d / DCAP64LVT
XXFILLER_259_1151 vdd_d vss_d / DCAP64LVT
XXFILLER_259_1587 vdd_d vss_d / DCAP64LVT
XXFILLER_259_1651 vdd_d vss_d / DCAP64LVT
XXFILLER_259_2087 vdd_d vss_d / DCAP64LVT
XXFILLER_259_2151 vdd_d vss_d / DCAP64LVT
XXFILLER_259_2215 vdd_d vss_d / DCAP64LVT
XXFILLER_259_2279 vdd_d vss_d / DCAP64LVT
XXplace2496 spi_bits[59] vdd_d vss_d net2496 / BUFFD6LVT
XXplace2498 spi_bits[58] vdd_d vss_d net2498 / BUFFD6LVT
XXplace2499 spi_bits[58] vdd_d vss_d net2499 / BUFFD6LVT
XXplace2501 spi_bits[57] vdd_d vss_d net2501 / BUFFD6LVT
XXplace2500 spi_bits[57] vdd_d vss_d net2500 / BUFFD6LVT
XXplace2503 spi_bits[56] vdd_d vss_d net2503 / BUFFD6LVT
XXplace2502 spi_bits[56] vdd_d vss_d net2502 / BUFFD6LVT
XXplace2504 spi_bits[55] vdd_d vss_d net2504 / BUFFD6LVT
XXplace2505 spi_bits[55] vdd_d vss_d net2505 / BUFFD6LVT
XXplace2506 spi_bits[54] vdd_d vss_d net2506 / BUFFD6LVT
XXplace2507 spi_bits[54] vdd_d vss_d net2507 / BUFFD6LVT
XXplace2508 spi_bits[53] vdd_d vss_d net2508 / BUFFD6LVT
XXplace2509 spi_bits[53] vdd_d vss_d net2509 / BUFFD6LVT
XXplace2510 spi_bits[52] vdd_d vss_d net2510 / BUFFD6LVT
XXplace2511 spi_bits[52] vdd_d vss_d net2511 / BUFFD6LVT
XXplace2512 spi_bits[51] vdd_d vss_d net2512 / BUFFD6LVT
XXplace2513 spi_bits[51] vdd_d vss_d net2513 / BUFFD6LVT
XXplace2514 spi_bits[50] vdd_d vss_d net2514 / BUFFD6LVT
XXplace2515 spi_bits[50] vdd_d vss_d net2515 / BUFFD6LVT
XXplace2517 net2516 vdd_d vss_d net2517 / BUFFD6LVT
XXplace2519 spi_bits[49] vdd_d vss_d net2519 / BUFFD6LVT
XXplace2520 spi_bits[49] vdd_d vss_d net2520 / BUFFD6LVT
XXplace2521 spi_bits[48] vdd_d vss_d net2521 / BUFFD6LVT
XXplace2522 spi_bits[48] vdd_d vss_d net2522 / BUFFD6LVT
XXplace2524 spi_bits[46] vdd_d vss_d net2524 / BUFFD6LVT
XXplace2525 spi_bits[46] vdd_d vss_d net2525 / BUFFD6LVT
XXplace2526 spi_bits[45] vdd_d vss_d net2526 / BUFFD6LVT
XXplace2527 spi_bits[45] vdd_d vss_d net2527 / BUFFD6LVT
XXplace2528 spi_bits[44] vdd_d vss_d net2528 / BUFFD6LVT
XXplace2529 spi_bits[44] vdd_d vss_d net2529 / BUFFD6LVT
XXplace2530 spi_bits[43] vdd_d vss_d net2530 / BUFFD6LVT
XXplace2531 spi_bits[43] vdd_d vss_d net2531 / BUFFD6LVT
XXplace2535 spi_bits[40] vdd_d vss_d net2535 / BUFFD6LVT
XXplace2534 spi_bits[40] vdd_d vss_d net2534 / BUFFD6LVT
XXplace2540 spi_bits[38] vdd_d vss_d net2540 / BUFFD6LVT
XXplace2541 spi_bits[38] vdd_d vss_d net2541 / BUFFD6LVT
XXplace2545 spi_bits[34] vdd_d vss_d net2545 / BUFFD6LVT
XXplace2546 spi_bits[34] vdd_d vss_d net2546 / BUFFD6LVT
XXplace2552 spi_bits[2] vdd_d vss_d net2552 / BUFFD6LVT
XXplace2551 spi_bits[30] vdd_d vss_d net2551 / BUFFD6LVT
XXplace2553 spi_bits[2] vdd_d vss_d net2553 / BUFFD6LVT
XXplace2550 spi_bits[30] vdd_d vss_d net2550 / BUFFD6LVT
XXplace2554 spi_bits[29] vdd_d vss_d net2554 / BUFFD6LVT
XXplace2555 spi_bits[29] vdd_d vss_d net2555 / BUFFD6LVT
XXplace2559 spi_bits[26] vdd_d vss_d net2559 / BUFFD6LVT
XXplace2558 spi_bits[26] vdd_d vss_d net2558 / BUFFD6LVT
XXplace2563 spi_bits[24] vdd_d vss_d net2563 / BUFFD6LVT
XXplace2561 spi_bits[25] vdd_d vss_d net2561 / BUFFD6LVT
XXplace2560 spi_bits[25] vdd_d vss_d net2560 / BUFFD6LVT
XXplace2562 spi_bits[24] vdd_d vss_d net2562 / BUFFD6LVT
XXplace2564 spi_bits[23] vdd_d vss_d net2564 / BUFFD6LVT
XXplace2565 spi_bits[23] vdd_d vss_d net2565 / BUFFD6LVT
XXplace2566 spi_bits[22] vdd_d vss_d net2566 / BUFFD6LVT
XXplace2567 spi_bits[22] vdd_d vss_d net2567 / BUFFD6LVT
XXplace2568 spi_bits[21] vdd_d vss_d net2568 / BUFFD6LVT
XXplace2569 spi_bits[21] vdd_d vss_d net2569 / BUFFD6LVT
XXplace2570 spi_bits[20] vdd_d vss_d net2570 / BUFFD6LVT
XXplace2571 spi_bits[20] vdd_d vss_d net2571 / BUFFD6LVT
XXplace2576 spi_bits[18] vdd_d vss_d net2576 / BUFFD6LVT
XXplace2573 spi_bits[19] vdd_d vss_d net2573 / BUFFD6LVT
XXplace2574 spi_bits[19] vdd_d vss_d net2574 / BUFFD6LVT
XXplace2575 spi_bits[18] vdd_d vss_d net2575 / BUFFD6LVT
XXplace2577 spi_bits[17] vdd_d vss_d net2577 / BUFFD6LVT
XXplace2578 spi_bits[17] vdd_d vss_d net2578 / BUFFD6LVT
XXplace2596 net2595 vdd_d vss_d net2596 / BUFFD6LVT
XXplace2593 net2592 vdd_d vss_d net2593 / BUFFD6LVT
XXplace2595 net2594 vdd_d vss_d net2595 / BUFFD6LVT
XXplace2594 net2593 vdd_d vss_d net2594 / BUFFD6LVT
XXplace2630 spi_bits[120] vdd_d vss_d net2630 / BUFFD6LVT
XXplace2583 spi_bits[175] vdd_d vss_d net2583 / BUFFD6LVT
XXplace2584 net2583 vdd_d vss_d net2584 / BUFFD6LVT
XXplace2587 spi_bits[16] vdd_d vss_d net2587 / BUFFD6LVT
XXplace2592 spi_bits[148] vdd_d vss_d net2592 / BUFFD6LVT
XXplace2696 net2695 vdd_d vss_d net2696 / BUFFD6LVT
XXplace2726 net2783 vdd_d vss_d net2726 / BUFFD6LVT
XXplace2497 spi_bits[59] vdd_d vss_d net2497 / BUFFD6LVT
XXplace2665 net2664 vdd_d vss_d net2665 / BUFFD6LVT
XXplace2632 spi_bits[11] vdd_d vss_d net2632 / BUFFD6LVT
XXplace2633 spi_bits[11] vdd_d vss_d net2633 / BUFFD6LVT
XXplace2537 net2536 vdd_d vss_d net2537 / BUFFD6LVT
XXplace2746 net2888 vdd_d vss_d net2746 / BUFFD6LVT
XXplace2750 net2887 vdd_d vss_d net2750 / BUFFD6LVT
XXplace2753 net2886 vdd_d vss_d net2753 / BUFFD6LVT
XXplace2757 net2802 vdd_d vss_d net2757 / BUFFD6LVT
XXplace2760 net2804 vdd_d vss_d net2760 / BUFFD6LVT
XXplace2493 spi_bits[60] vdd_d vss_d net2493 / BUFFD6LVT
XXplace2494 spi_bits[60] vdd_d vss_d net2494 / BUFFD6LVT
XXplace2491 spi_bits[61] vdd_d vss_d net2491 / BUFFD6LVT
XXplace2492 spi_bits[61] vdd_d vss_d net2492 / BUFFD6LVT
XXplace2488 net2487 vdd_d vss_d net2488 / BUFFD6LVT
XXplace2486 spi_bits[6] vdd_d vss_d net2486 / BUFFD6LVT
XXplace2485 spi_bits[6] vdd_d vss_d net2485 / BUFFD6LVT
XXplace2482 spi_bits[7] vdd_d vss_d net2482 / BUFFD6LVT
XXplace2483 spi_bits[7] vdd_d vss_d net2483 / BUFFD6LVT
XXplace2477 net2772 vdd_d vss_d net2477 / BUFFD6LVT
XXplace2588 spi_bits[16] vdd_d vss_d net2588 / BUFFD6LVT
XXplace2622 spi_bits[127] vdd_d vss_d net2622 / BUFFD6LVT
XXplace2729 net2890 vdd_d vss_d net2729 / BUFFD6LVT
XXplace2730 net2729 vdd_d vss_d net2730 / BUFFD6LVT
XXplace2739 net2895 vdd_d vss_d net2739 / BUFFD6LVT
XXplace2742 net2790 vdd_d vss_d net2742 / BUFFD6LVT
XXplace2743 net2742 vdd_d vss_d net2743 / BUFFD6LVT
XXplace2747 net2746 vdd_d vss_d net2747 / BUFFD6LVT
XXplace2754 net2753 vdd_d vss_d net2754 / BUFFD6LVT
XXplace2481 spi_bits[8] vdd_d vss_d net2481 / CKBD16LVT
XXplace2523 spi_bits[47] vdd_d vss_d net2523 / CKBD16LVT
XXplace2532 spi_bits[42] vdd_d vss_d net2532 / CKBD16LVT
XXplace2533 spi_bits[41] vdd_d vss_d net2533 / CKBD16LVT
XXplace2539 spi_bits[39] vdd_d vss_d net2539 / CKBD16LVT
XXplace2542 spi_bits[37] vdd_d vss_d net2542 / CKBD16LVT
XXplace2543 spi_bits[36] vdd_d vss_d net2543 / CKBD16LVT
XXplace2544 spi_bits[35] vdd_d vss_d net2544 / CKBD16LVT
XXplace2547 spi_bits[33] vdd_d vss_d net2547 / CKBD16LVT
XXplace2548 spi_bits[32] vdd_d vss_d net2548 / CKBD16LVT
XXplace2549 spi_bits[31] vdd_d vss_d net2549 / CKBD16LVT
XXplace2556 spi_bits[28] vdd_d vss_d net2556 / CKBD16LVT
XXplace2557 spi_bits[27] vdd_d vss_d net2557 / CKBD16LVT
XXplace2572 spi_bits[1] vdd_d vss_d net2572 / CKBD16LVT
XXplace2589 spi_bits[15] vdd_d vss_d net2589 / CKBD16LVT
XXplace2591 spi_bits[14] vdd_d vss_d net2591 / CKBD16LVT
XXplace2646 spi_bits[10] vdd_d vss_d net2646 / CKBD16LVT
XXplace2657 spi_bits[0] vdd_d vss_d net2657 / CKBD16LVT
XXplace2469 spi_bits[9] vdd_d vss_d net2469 / CKBD16LVT
XXplace2495 spi_bits[5] vdd_d vss_d net2495 / CKBD16LVT
XXplace2490 spi_bits[62] vdd_d vss_d net2490 / CKBD16LVT
XXplace2608 spi_bits[13] vdd_d vss_d net2608 / CKBD16LVT
XXplace2619 spi_bits[12] vdd_d vss_d net2619 / CKBD16LVT
XXFILLER_19_1162 vdd_d vss_d / DCAP4LVT
XXFILLER_15_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_14_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_13_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_12_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_10_1249 vdd_d vss_d / DCAP4LVT
XXFILLER_10_856 vdd_d vss_d / DCAP4LVT
XXFILLER_9_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_7_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_10_816 vdd_d vss_d / DCAP4LVT
XXFILLER_6_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_8_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_5_749 vdd_d vss_d / DCAP4LVT
XXFILLER_4_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_4_402 vdd_d vss_d / DCAP4LVT
XXFILLER_3_384 vdd_d vss_d / DCAP4LVT
XXFILLER_2_2346 vdd_d vss_d / DCAP4LVT
XXFILLER_2_777 vdd_d vss_d / DCAP4LVT
XXFILLER_2_749 vdd_d vss_d / DCAP4LVT
XXFILLER_2_448 vdd_d vss_d / DCAP4LVT
XXFILLER_2_812 vdd_d vss_d / DCAP4LVT
XXFILLER_2_615 vdd_d vss_d / DCAP4LVT
XXFILLER_1_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_16_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_17_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_18_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_19_536 vdd_d vss_d / DCAP4LVT
XXFILLER_0_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_20_1159 vdd_d vss_d / DCAP4LVT
XXFILLER_20_1204 vdd_d vss_d / DCAP4LVT
XXFILLER_20_1612 vdd_d vss_d / DCAP4LVT
XXFILLER_20_1716 vdd_d vss_d / DCAP4LVT
XXFILLER_20_2346 vdd_d vss_d / DCAP4LVT
XXFILLER_21_1224 vdd_d vss_d / DCAP4LVT
XXFILLER_21_1605 vdd_d vss_d / DCAP4LVT
XXFILLER_22_1120 vdd_d vss_d / DCAP4LVT
XXFILLER_22_1138 vdd_d vss_d / DCAP4LVT
XXFILLER_22_1232 vdd_d vss_d / DCAP4LVT
XXFILLER_22_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_23_449 vdd_d vss_d / DCAP4LVT
XXFILLER_23_1157 vdd_d vss_d / DCAP4LVT
XXFILLER_23_1194 vdd_d vss_d / DCAP4LVT
XXFILLER_23_1226 vdd_d vss_d / DCAP4LVT
XXFILLER_23_1347 vdd_d vss_d / DCAP4LVT
XXFILLER_23_2345 vdd_d vss_d / DCAP4LVT
XXFILLER_24_400 vdd_d vss_d / DCAP4LVT
XXFILLER_24_441 vdd_d vss_d / DCAP4LVT
XXFILLER_24_1067 vdd_d vss_d / DCAP4LVT
XXFILLER_25_1117 vdd_d vss_d / DCAP4LVT
XXFILLER_25_1225 vdd_d vss_d / DCAP4LVT
XXFILLER_25_1236 vdd_d vss_d / DCAP4LVT
XXFILLER_25_2346 vdd_d vss_d / DCAP4LVT
XXFILLER_26_392 vdd_d vss_d / DCAP4LVT
XXFILLER_26_442 vdd_d vss_d / DCAP4LVT
XXFILLER_26_1043 vdd_d vss_d / DCAP4LVT
XXFILLER_26_1069 vdd_d vss_d / DCAP4LVT
XXFILLER_26_1731 vdd_d vss_d / DCAP4LVT
XXFILLER_27_400 vdd_d vss_d / DCAP4LVT
XXFILLER_27_440 vdd_d vss_d / DCAP4LVT
XXFILLER_27_450 vdd_d vss_d / DCAP4LVT
XXFILLER_27_1032 vdd_d vss_d / DCAP4LVT
XXFILLER_27_1042 vdd_d vss_d / DCAP4LVT
XXFILLER_27_1062 vdd_d vss_d / DCAP4LVT
XXFILLER_27_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_28_449 vdd_d vss_d / DCAP4LVT
XXFILLER_28_593 vdd_d vss_d / DCAP4LVT
XXFILLER_28_1144 vdd_d vss_d / DCAP4LVT
XXFILLER_28_2345 vdd_d vss_d / DCAP4LVT
XXFILLER_29_440 vdd_d vss_d / DCAP4LVT
XXFILLER_29_897 vdd_d vss_d / DCAP4LVT
XXFILLER_29_1333 vdd_d vss_d / DCAP4LVT
XXFILLER_29_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_30_994 vdd_d vss_d / DCAP4LVT
XXFILLER_30_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_31_499 vdd_d vss_d / DCAP4LVT
XXFILLER_31_782 vdd_d vss_d / DCAP4LVT
XXFILLER_31_1464 vdd_d vss_d / DCAP4LVT
XXFILLER_31_1872 vdd_d vss_d / DCAP4LVT
XXFILLER_31_1882 vdd_d vss_d / DCAP4LVT
XXFILLER_32_788 vdd_d vss_d / DCAP4LVT
XXFILLER_32_982 vdd_d vss_d / DCAP4LVT
XXFILLER_32_1393 vdd_d vss_d / DCAP4LVT
XXFILLER_32_1419 vdd_d vss_d / DCAP4LVT
XXFILLER_32_1469 vdd_d vss_d / DCAP4LVT
XXFILLER_33_416 vdd_d vss_d / DCAP4LVT
XXFILLER_33_926 vdd_d vss_d / DCAP4LVT
XXFILLER_33_1184 vdd_d vss_d / DCAP4LVT
XXFILLER_33_1453 vdd_d vss_d / DCAP4LVT
XXFILLER_33_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_34_996 vdd_d vss_d / DCAP4LVT
XXFILLER_34_1091 vdd_d vss_d / DCAP4LVT
XXFILLER_34_1138 vdd_d vss_d / DCAP4LVT
XXFILLER_34_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_35_480 vdd_d vss_d / DCAP4LVT
XXFILLER_35_507 vdd_d vss_d / DCAP4LVT
XXFILLER_35_523 vdd_d vss_d / DCAP4LVT
XXFILLER_35_580 vdd_d vss_d / DCAP4LVT
XXFILLER_35_948 vdd_d vss_d / DCAP4LVT
XXFILLER_35_1160 vdd_d vss_d / DCAP4LVT
XXFILLER_35_1299 vdd_d vss_d / DCAP4LVT
XXFILLER_35_1421 vdd_d vss_d / DCAP4LVT
XXFILLER_35_1433 vdd_d vss_d / DCAP4LVT
XXFILLER_35_1480 vdd_d vss_d / DCAP4LVT
XXFILLER_35_1492 vdd_d vss_d / DCAP4LVT
XXFILLER_36_408 vdd_d vss_d / DCAP4LVT
XXFILLER_36_858 vdd_d vss_d / DCAP4LVT
XXFILLER_36_897 vdd_d vss_d / DCAP4LVT
XXFILLER_36_948 vdd_d vss_d / DCAP4LVT
XXFILLER_36_1113 vdd_d vss_d / DCAP4LVT
XXFILLER_36_1260 vdd_d vss_d / DCAP4LVT
XXFILLER_36_1280 vdd_d vss_d / DCAP4LVT
XXFILLER_36_1290 vdd_d vss_d / DCAP4LVT
XXFILLER_36_1404 vdd_d vss_d / DCAP4LVT
XXFILLER_36_1424 vdd_d vss_d / DCAP4LVT
XXFILLER_36_1880 vdd_d vss_d / DCAP4LVT
XXFILLER_37_384 vdd_d vss_d / DCAP4LVT
XXFILLER_37_477 vdd_d vss_d / DCAP4LVT
XXFILLER_37_533 vdd_d vss_d / DCAP4LVT
XXFILLER_37_829 vdd_d vss_d / DCAP4LVT
XXFILLER_37_893 vdd_d vss_d / DCAP4LVT
XXFILLER_37_934 vdd_d vss_d / DCAP4LVT
XXFILLER_37_1457 vdd_d vss_d / DCAP4LVT
XXFILLER_37_1634 vdd_d vss_d / DCAP4LVT
XXFILLER_37_1828 vdd_d vss_d / DCAP4LVT
XXFILLER_37_1912 vdd_d vss_d / DCAP4LVT
XXFILLER_38_637 vdd_d vss_d / DCAP4LVT
XXFILLER_38_808 vdd_d vss_d / DCAP4LVT
XXFILLER_38_865 vdd_d vss_d / DCAP4LVT
XXFILLER_38_1197 vdd_d vss_d / DCAP4LVT
XXFILLER_38_1353 vdd_d vss_d / DCAP4LVT
XXFILLER_38_1451 vdd_d vss_d / DCAP4LVT
XXFILLER_38_1507 vdd_d vss_d / DCAP4LVT
XXFILLER_38_1591 vdd_d vss_d / DCAP4LVT
XXFILLER_38_1630 vdd_d vss_d / DCAP4LVT
XXFILLER_38_1845 vdd_d vss_d / DCAP4LVT
XXFILLER_38_2346 vdd_d vss_d / DCAP4LVT
XXFILLER_39_384 vdd_d vss_d / DCAP4LVT
XXFILLER_39_425 vdd_d vss_d / DCAP4LVT
XXFILLER_39_752 vdd_d vss_d / DCAP4LVT
XXFILLER_39_895 vdd_d vss_d / DCAP4LVT
XXFILLER_39_949 vdd_d vss_d / DCAP4LVT
XXFILLER_39_1192 vdd_d vss_d / DCAP4LVT
XXFILLER_39_1243 vdd_d vss_d / DCAP4LVT
XXFILLER_39_1378 vdd_d vss_d / DCAP4LVT
XXFILLER_39_1478 vdd_d vss_d / DCAP4LVT
XXFILLER_39_1533 vdd_d vss_d / DCAP4LVT
XXFILLER_39_1859 vdd_d vss_d / DCAP4LVT
XXFILLER_39_1936 vdd_d vss_d / DCAP4LVT
XXFILLER_39_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_40_384 vdd_d vss_d / DCAP4LVT
XXFILLER_40_433 vdd_d vss_d / DCAP4LVT
XXFILLER_40_541 vdd_d vss_d / DCAP4LVT
XXFILLER_40_768 vdd_d vss_d / DCAP4LVT
XXFILLER_40_974 vdd_d vss_d / DCAP4LVT
XXFILLER_40_984 vdd_d vss_d / DCAP4LVT
XXFILLER_40_1019 vdd_d vss_d / DCAP4LVT
XXFILLER_40_1054 vdd_d vss_d / DCAP4LVT
XXFILLER_40_1112 vdd_d vss_d / DCAP4LVT
XXFILLER_40_1267 vdd_d vss_d / DCAP4LVT
XXFILLER_40_1600 vdd_d vss_d / DCAP4LVT
XXFILLER_40_1850 vdd_d vss_d / DCAP4LVT
XXFILLER_41_438 vdd_d vss_d / DCAP4LVT
XXFILLER_41_846 vdd_d vss_d / DCAP4LVT
XXFILLER_41_953 vdd_d vss_d / DCAP4LVT
XXFILLER_41_1044 vdd_d vss_d / DCAP4LVT
XXFILLER_41_1220 vdd_d vss_d / DCAP4LVT
XXFILLER_41_1500 vdd_d vss_d / DCAP4LVT
XXFILLER_41_1803 vdd_d vss_d / DCAP4LVT
XXFILLER_41_1819 vdd_d vss_d / DCAP4LVT
XXFILLER_41_1867 vdd_d vss_d / DCAP4LVT
XXFILLER_41_1908 vdd_d vss_d / DCAP4LVT
XXFILLER_41_1948 vdd_d vss_d / DCAP4LVT
XXFILLER_42_755 vdd_d vss_d / DCAP4LVT
XXFILLER_42_821 vdd_d vss_d / DCAP4LVT
XXFILLER_42_860 vdd_d vss_d / DCAP4LVT
XXFILLER_42_878 vdd_d vss_d / DCAP4LVT
XXFILLER_42_920 vdd_d vss_d / DCAP4LVT
XXFILLER_42_983 vdd_d vss_d / DCAP4LVT
XXFILLER_42_1119 vdd_d vss_d / DCAP4LVT
XXFILLER_42_1244 vdd_d vss_d / DCAP4LVT
XXFILLER_42_1327 vdd_d vss_d / DCAP4LVT
XXFILLER_42_1363 vdd_d vss_d / DCAP4LVT
XXFILLER_42_1375 vdd_d vss_d / DCAP4LVT
XXFILLER_42_1475 vdd_d vss_d / DCAP4LVT
XXFILLER_42_1511 vdd_d vss_d / DCAP4LVT
XXFILLER_42_1561 vdd_d vss_d / DCAP4LVT
XXFILLER_42_1605 vdd_d vss_d / DCAP4LVT
XXFILLER_42_1663 vdd_d vss_d / DCAP4LVT
XXFILLER_42_1883 vdd_d vss_d / DCAP4LVT
XXFILLER_42_1914 vdd_d vss_d / DCAP4LVT
XXFILLER_42_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_43_384 vdd_d vss_d / DCAP4LVT
XXFILLER_43_707 vdd_d vss_d / DCAP4LVT
XXFILLER_43_740 vdd_d vss_d / DCAP4LVT
XXFILLER_43_895 vdd_d vss_d / DCAP4LVT
XXFILLER_43_1084 vdd_d vss_d / DCAP4LVT
XXFILLER_43_1148 vdd_d vss_d / DCAP4LVT
XXFILLER_43_1206 vdd_d vss_d / DCAP4LVT
XXFILLER_43_1233 vdd_d vss_d / DCAP4LVT
XXFILLER_43_1365 vdd_d vss_d / DCAP4LVT
XXFILLER_43_1439 vdd_d vss_d / DCAP4LVT
XXFILLER_43_1491 vdd_d vss_d / DCAP4LVT
XXFILLER_43_1647 vdd_d vss_d / DCAP4LVT
XXFILLER_43_1801 vdd_d vss_d / DCAP4LVT
XXFILLER_43_1886 vdd_d vss_d / DCAP4LVT
XXFILLER_43_2346 vdd_d vss_d / DCAP4LVT
XXFILLER_44_383 vdd_d vss_d / DCAP4LVT
XXFILLER_44_424 vdd_d vss_d / DCAP4LVT
XXFILLER_44_444 vdd_d vss_d / DCAP4LVT
XXFILLER_44_469 vdd_d vss_d / DCAP4LVT
XXFILLER_44_481 vdd_d vss_d / DCAP4LVT
XXFILLER_44_810 vdd_d vss_d / DCAP4LVT
XXFILLER_44_826 vdd_d vss_d / DCAP4LVT
XXFILLER_44_912 vdd_d vss_d / DCAP4LVT
XXFILLER_44_1002 vdd_d vss_d / DCAP4LVT
XXFILLER_44_1083 vdd_d vss_d / DCAP4LVT
XXFILLER_44_1126 vdd_d vss_d / DCAP4LVT
XXFILLER_44_1151 vdd_d vss_d / DCAP4LVT
XXFILLER_44_1219 vdd_d vss_d / DCAP4LVT
XXFILLER_44_1267 vdd_d vss_d / DCAP4LVT
XXFILLER_44_1369 vdd_d vss_d / DCAP4LVT
XXFILLER_44_1477 vdd_d vss_d / DCAP4LVT
XXFILLER_44_1533 vdd_d vss_d / DCAP4LVT
XXFILLER_44_1833 vdd_d vss_d / DCAP4LVT
XXFILLER_44_1887 vdd_d vss_d / DCAP4LVT
XXFILLER_44_1898 vdd_d vss_d / DCAP4LVT
XXFILLER_44_1918 vdd_d vss_d / DCAP4LVT
XXFILLER_44_1936 vdd_d vss_d / DCAP4LVT
XXFILLER_44_2346 vdd_d vss_d / DCAP4LVT
XXFILLER_45_832 vdd_d vss_d / DCAP4LVT
XXFILLER_45_1589 vdd_d vss_d / DCAP4LVT
XXFILLER_46_1538 vdd_d vss_d / DCAP4LVT
XXFILLER_46_1688 vdd_d vss_d / DCAP4LVT
XXFILLER_46_1701 vdd_d vss_d / DCAP4LVT
XXFILLER_46_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_47_664 vdd_d vss_d / DCAP4LVT
XXFILLER_47_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_48_88 vdd_d vss_d / DCAP4LVT
XXFILLER_48_914 vdd_d vss_d / DCAP4LVT
XXFILLER_48_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_49_408 vdd_d vss_d / DCAP4LVT
XXFILLER_49_1487 vdd_d vss_d / DCAP4LVT
XXFILLER_49_2345 vdd_d vss_d / DCAP4LVT
XXFILLER_50_410 vdd_d vss_d / DCAP4LVT
XXFILLER_50_819 vdd_d vss_d / DCAP4LVT
XXFILLER_50_1485 vdd_d vss_d / DCAP4LVT
XXFILLER_50_1737 vdd_d vss_d / DCAP4LVT
XXFILLER_50_1914 vdd_d vss_d / DCAP4LVT
XXFILLER_52_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_53_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_54_901 vdd_d vss_d / DCAP4LVT
XXFILLER_54_1943 vdd_d vss_d / DCAP4LVT
XXFILLER_55_424 vdd_d vss_d / DCAP4LVT
XXFILLER_55_885 vdd_d vss_d / DCAP4LVT
XXFILLER_55_1944 vdd_d vss_d / DCAP4LVT
XXFILLER_55_2346 vdd_d vss_d / DCAP4LVT
XXFILLER_56_256 vdd_d vss_d / DCAP4LVT
XXFILLER_56_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_57_256 vdd_d vss_d / DCAP4LVT
XXFILLER_57_1667 vdd_d vss_d / DCAP4LVT
XXFILLER_57_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_58_256 vdd_d vss_d / DCAP4LVT
XXFILLER_58_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_59_256 vdd_d vss_d / DCAP4LVT
XXFILLER_59_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_60_256 vdd_d vss_d / DCAP4LVT
XXFILLER_60_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_61_256 vdd_d vss_d / DCAP4LVT
XXFILLER_61_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_62_256 vdd_d vss_d / DCAP4LVT
XXFILLER_62_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_63_256 vdd_d vss_d / DCAP4LVT
XXFILLER_63_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_64_256 vdd_d vss_d / DCAP4LVT
XXFILLER_64_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_65_256 vdd_d vss_d / DCAP4LVT
XXFILLER_65_755 vdd_d vss_d / DCAP4LVT
XXFILLER_65_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_66_256 vdd_d vss_d / DCAP4LVT
XXFILLER_66_723 vdd_d vss_d / DCAP4LVT
XXFILLER_66_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_67_256 vdd_d vss_d / DCAP4LVT
XXFILLER_67_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_68_256 vdd_d vss_d / DCAP4LVT
XXFILLER_68_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_69_240 vdd_d vss_d / DCAP4LVT
XXFILLER_69_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_70_256 vdd_d vss_d / DCAP4LVT
XXFILLER_70_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_71_256 vdd_d vss_d / DCAP4LVT
XXFILLER_71_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_72_256 vdd_d vss_d / DCAP4LVT
XXFILLER_72_1111 vdd_d vss_d / DCAP4LVT
XXFILLER_72_1256 vdd_d vss_d / DCAP4LVT
XXFILLER_72_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_73_248 vdd_d vss_d / DCAP4LVT
XXFILLER_73_2346 vdd_d vss_d / DCAP4LVT
XXFILLER_74_256 vdd_d vss_d / DCAP4LVT
XXFILLER_74_1127 vdd_d vss_d / DCAP4LVT
XXFILLER_74_1257 vdd_d vss_d / DCAP4LVT
XXFILLER_74_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_75_256 vdd_d vss_d / DCAP4LVT
XXFILLER_75_1747 vdd_d vss_d / DCAP4LVT
XXFILLER_75_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_76_248 vdd_d vss_d / DCAP4LVT
XXFILLER_76_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_77_256 vdd_d vss_d / DCAP4LVT
XXFILLER_77_1207 vdd_d vss_d / DCAP4LVT
XXFILLER_77_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_78_256 vdd_d vss_d / DCAP4LVT
XXFILLER_78_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_79_256 vdd_d vss_d / DCAP4LVT
XXFILLER_79_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_80_256 vdd_d vss_d / DCAP4LVT
XXFILLER_80_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_81_256 vdd_d vss_d / DCAP4LVT
XXFILLER_81_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_82_256 vdd_d vss_d / DCAP4LVT
XXFILLER_82_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_83_224 vdd_d vss_d / DCAP4LVT
XXFILLER_83_1239 vdd_d vss_d / DCAP4LVT
XXFILLER_83_1258 vdd_d vss_d / DCAP4LVT
XXFILLER_83_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_84_256 vdd_d vss_d / DCAP4LVT
XXFILLER_84_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_85_256 vdd_d vss_d / DCAP4LVT
XXFILLER_85_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_86_256 vdd_d vss_d / DCAP4LVT
XXFILLER_86_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_87_256 vdd_d vss_d / DCAP4LVT
XXFILLER_87_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_88_256 vdd_d vss_d / DCAP4LVT
XXFILLER_88_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_89_256 vdd_d vss_d / DCAP4LVT
XXFILLER_89_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_90_256 vdd_d vss_d / DCAP4LVT
XXFILLER_90_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_91_256 vdd_d vss_d / DCAP4LVT
XXFILLER_91_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_92_256 vdd_d vss_d / DCAP4LVT
XXFILLER_92_1223 vdd_d vss_d / DCAP4LVT
XXFILLER_92_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_93_256 vdd_d vss_d / DCAP4LVT
XXFILLER_93_1739 vdd_d vss_d / DCAP4LVT
XXFILLER_93_1759 vdd_d vss_d / DCAP4LVT
XXFILLER_93_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_94_256 vdd_d vss_d / DCAP4LVT
XXFILLER_94_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_95_408 vdd_d vss_d / DCAP4LVT
XXFILLER_95_447 vdd_d vss_d / DCAP4LVT
XXFILLER_95_964 vdd_d vss_d / DCAP4LVT
XXFILLER_95_1412 vdd_d vss_d / DCAP4LVT
XXFILLER_95_1438 vdd_d vss_d / DCAP4LVT
XXFILLER_96_360 vdd_d vss_d / DCAP4LVT
XXFILLER_97_1446 vdd_d vss_d / DCAP4LVT
XXFILLER_98_1617 vdd_d vss_d / DCAP4LVT
XXFILLER_99_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_100_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_102_672 vdd_d vss_d / DCAP4LVT
XXFILLER_103_1616 vdd_d vss_d / DCAP4LVT
XXFILLER_103_1908 vdd_d vss_d / DCAP4LVT
XXFILLER_104_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_105_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_106_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_107_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_109_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_110_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_111_1463 vdd_d vss_d / DCAP4LVT
XXFILLER_112_256 vdd_d vss_d / DCAP4LVT
XXFILLER_112_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_113_256 vdd_d vss_d / DCAP4LVT
XXFILLER_113_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_114_256 vdd_d vss_d / DCAP4LVT
XXFILLER_114_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_115_256 vdd_d vss_d / DCAP4LVT
XXFILLER_115_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_116_256 vdd_d vss_d / DCAP4LVT
XXFILLER_116_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_117_256 vdd_d vss_d / DCAP4LVT
XXFILLER_117_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_118_256 vdd_d vss_d / DCAP4LVT
XXFILLER_118_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_119_256 vdd_d vss_d / DCAP4LVT
XXFILLER_119_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_120_256 vdd_d vss_d / DCAP4LVT
XXFILLER_120_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_121_256 vdd_d vss_d / DCAP4LVT
XXFILLER_121_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_122_256 vdd_d vss_d / DCAP4LVT
XXFILLER_122_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_123_256 vdd_d vss_d / DCAP4LVT
XXFILLER_123_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_124_256 vdd_d vss_d / DCAP4LVT
XXFILLER_124_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_125_256 vdd_d vss_d / DCAP4LVT
XXFILLER_125_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_126_256 vdd_d vss_d / DCAP4LVT
XXFILLER_126_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_127_256 vdd_d vss_d / DCAP4LVT
XXFILLER_127_1747 vdd_d vss_d / DCAP4LVT
XXFILLER_127_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_128_256 vdd_d vss_d / DCAP4LVT
XXFILLER_128_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_129_256 vdd_d vss_d / DCAP4LVT
XXFILLER_129_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_130_256 vdd_d vss_d / DCAP4LVT
XXFILLER_130_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_132_256 vdd_d vss_d / DCAP4LVT
XXFILLER_132_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_133_256 vdd_d vss_d / DCAP4LVT
XXFILLER_133_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_134_256 vdd_d vss_d / DCAP4LVT
XXFILLER_134_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_135_256 vdd_d vss_d / DCAP4LVT
XXFILLER_135_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_136_256 vdd_d vss_d / DCAP4LVT
XXFILLER_136_756 vdd_d vss_d / DCAP4LVT
XXFILLER_136_1757 vdd_d vss_d / DCAP4LVT
XXFILLER_136_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_137_256 vdd_d vss_d / DCAP4LVT
XXFILLER_137_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_138_256 vdd_d vss_d / DCAP4LVT
XXFILLER_138_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_139_256 vdd_d vss_d / DCAP4LVT
XXFILLER_139_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_140_256 vdd_d vss_d / DCAP4LVT
XXFILLER_140_1175 vdd_d vss_d / DCAP4LVT
XXFILLER_140_1256 vdd_d vss_d / DCAP4LVT
XXFILLER_140_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_141_256 vdd_d vss_d / DCAP4LVT
XXFILLER_141_1151 vdd_d vss_d / DCAP4LVT
XXFILLER_141_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_142_256 vdd_d vss_d / DCAP4LVT
XXFILLER_142_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_143_256 vdd_d vss_d / DCAP4LVT
XXFILLER_143_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_144_256 vdd_d vss_d / DCAP4LVT
XXFILLER_144_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_145_256 vdd_d vss_d / DCAP4LVT
XXFILLER_145_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_146_256 vdd_d vss_d / DCAP4LVT
XXFILLER_146_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_147_256 vdd_d vss_d / DCAP4LVT
XXFILLER_147_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_148_256 vdd_d vss_d / DCAP4LVT
XXFILLER_148_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_149_256 vdd_d vss_d / DCAP4LVT
XXFILLER_149_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_150_432 vdd_d vss_d / DCAP4LVT
XXFILLER_150_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_151_440 vdd_d vss_d / DCAP4LVT
XXFILLER_151_1415 vdd_d vss_d / DCAP4LVT
XXFILLER_152_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_153_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_154_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_155_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_156_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_157_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_158_688 vdd_d vss_d / DCAP4LVT
XXFILLER_158_2346 vdd_d vss_d / DCAP4LVT
XXFILLER_159_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_160_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_161_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_162_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_163_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_164_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_165_1864 vdd_d vss_d / DCAP4LVT
XXFILLER_165_2345 vdd_d vss_d / DCAP4LVT
XXFILLER_166_1859 vdd_d vss_d / DCAP4LVT
XXFILLER_167_256 vdd_d vss_d / DCAP4LVT
XXFILLER_167_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_168_256 vdd_d vss_d / DCAP4LVT
XXFILLER_168_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_169_256 vdd_d vss_d / DCAP4LVT
XXFILLER_169_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_170_256 vdd_d vss_d / DCAP4LVT
XXFILLER_170_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_171_256 vdd_d vss_d / DCAP4LVT
XXFILLER_171_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_172_256 vdd_d vss_d / DCAP4LVT
XXFILLER_172_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_173_256 vdd_d vss_d / DCAP4LVT
XXFILLER_173_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_174_256 vdd_d vss_d / DCAP4LVT
XXFILLER_174_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_175_256 vdd_d vss_d / DCAP4LVT
XXFILLER_175_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_176_256 vdd_d vss_d / DCAP4LVT
XXFILLER_176_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_177_256 vdd_d vss_d / DCAP4LVT
XXFILLER_177_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_178_256 vdd_d vss_d / DCAP4LVT
XXFILLER_178_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_179_256 vdd_d vss_d / DCAP4LVT
XXFILLER_179_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_180_256 vdd_d vss_d / DCAP4LVT
XXFILLER_180_1175 vdd_d vss_d / DCAP4LVT
XXFILLER_180_1256 vdd_d vss_d / DCAP4LVT
XXFILLER_180_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_181_256 vdd_d vss_d / DCAP4LVT
XXFILLER_181_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_182_256 vdd_d vss_d / DCAP4LVT
XXFILLER_182_1238 vdd_d vss_d / DCAP4LVT
XXFILLER_182_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_183_256 vdd_d vss_d / DCAP4LVT
XXFILLER_183_1248 vdd_d vss_d / DCAP4LVT
XXFILLER_183_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_184_256 vdd_d vss_d / DCAP4LVT
XXFILLER_184_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_185_256 vdd_d vss_d / DCAP4LVT
XXFILLER_185_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_186_256 vdd_d vss_d / DCAP4LVT
XXFILLER_186_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_187_256 vdd_d vss_d / DCAP4LVT
XXFILLER_187_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_188_256 vdd_d vss_d / DCAP4LVT
XXFILLER_188_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_189_256 vdd_d vss_d / DCAP4LVT
XXFILLER_189_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_190_256 vdd_d vss_d / DCAP4LVT
XXFILLER_190_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_191_256 vdd_d vss_d / DCAP4LVT
XXFILLER_191_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_192_256 vdd_d vss_d / DCAP4LVT
XXFILLER_192_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_193_256 vdd_d vss_d / DCAP4LVT
XXFILLER_193_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_194_256 vdd_d vss_d / DCAP4LVT
XXFILLER_194_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_195_256 vdd_d vss_d / DCAP4LVT
XXFILLER_195_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_196_256 vdd_d vss_d / DCAP4LVT
XXFILLER_196_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_197_256 vdd_d vss_d / DCAP4LVT
XXFILLER_197_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_198_256 vdd_d vss_d / DCAP4LVT
XXFILLER_198_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_199_256 vdd_d vss_d / DCAP4LVT
XXFILLER_199_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_200_256 vdd_d vss_d / DCAP4LVT
XXFILLER_200_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_201_256 vdd_d vss_d / DCAP4LVT
XXFILLER_201_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_202_256 vdd_d vss_d / DCAP4LVT
XXFILLER_202_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_203_256 vdd_d vss_d / DCAP4LVT
XXFILLER_203_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_204_256 vdd_d vss_d / DCAP4LVT
XXFILLER_204_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_205_256 vdd_d vss_d / DCAP4LVT
XXFILLER_205_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_206_432 vdd_d vss_d / DCAP4LVT
XXFILLER_206_943 vdd_d vss_d / DCAP4LVT
XXFILLER_206_1428 vdd_d vss_d / DCAP4LVT
XXFILLER_207_936 vdd_d vss_d / DCAP4LVT
XXFILLER_208_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_209_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_210_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_211_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_212_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_213_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_214_696 vdd_d vss_d / DCAP4LVT
XXFILLER_214_1925 vdd_d vss_d / DCAP4LVT
XXFILLER_214_2345 vdd_d vss_d / DCAP4LVT
XXFILLER_215_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_216_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_217_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_218_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_219_904 vdd_d vss_d / DCAP4LVT
XXFILLER_219_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_220_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_221_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_222_2344 vdd_d vss_d / DCAP4LVT
XXFILLER_223_256 vdd_d vss_d / DCAP4LVT
XXFILLER_223_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_224_256 vdd_d vss_d / DCAP4LVT
XXFILLER_224_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_225_256 vdd_d vss_d / DCAP4LVT
XXFILLER_225_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_226_256 vdd_d vss_d / DCAP4LVT
XXFILLER_226_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_227_256 vdd_d vss_d / DCAP4LVT
XXFILLER_227_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_228_256 vdd_d vss_d / DCAP4LVT
XXFILLER_228_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_229_256 vdd_d vss_d / DCAP4LVT
XXFILLER_229_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_230_256 vdd_d vss_d / DCAP4LVT
XXFILLER_230_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_231_256 vdd_d vss_d / DCAP4LVT
XXFILLER_231_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_232_256 vdd_d vss_d / DCAP4LVT
XXFILLER_232_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_233_256 vdd_d vss_d / DCAP4LVT
XXFILLER_233_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_234_256 vdd_d vss_d / DCAP4LVT
XXFILLER_234_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_235_256 vdd_d vss_d / DCAP4LVT
XXFILLER_235_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_236_256 vdd_d vss_d / DCAP4LVT
XXFILLER_236_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_237_256 vdd_d vss_d / DCAP4LVT
XXFILLER_237_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_238_256 vdd_d vss_d / DCAP4LVT
XXFILLER_238_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_239_256 vdd_d vss_d / DCAP4LVT
XXFILLER_239_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_240_256 vdd_d vss_d / DCAP4LVT
XXFILLER_240_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_241_256 vdd_d vss_d / DCAP4LVT
XXFILLER_241_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_242_256 vdd_d vss_d / DCAP4LVT
XXFILLER_242_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_243_256 vdd_d vss_d / DCAP4LVT
XXFILLER_243_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_244_256 vdd_d vss_d / DCAP4LVT
XXFILLER_244_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_245_256 vdd_d vss_d / DCAP4LVT
XXFILLER_245_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_246_256 vdd_d vss_d / DCAP4LVT
XXFILLER_246_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_247_256 vdd_d vss_d / DCAP4LVT
XXFILLER_247_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_248_256 vdd_d vss_d / DCAP4LVT
XXFILLER_248_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_249_256 vdd_d vss_d / DCAP4LVT
XXFILLER_249_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_250_256 vdd_d vss_d / DCAP4LVT
XXFILLER_250_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_251_256 vdd_d vss_d / DCAP4LVT
XXFILLER_251_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_252_256 vdd_d vss_d / DCAP4LVT
XXFILLER_252_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_253_256 vdd_d vss_d / DCAP4LVT
XXFILLER_253_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_254_256 vdd_d vss_d / DCAP4LVT
XXFILLER_254_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_255_256 vdd_d vss_d / DCAP4LVT
XXFILLER_255_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_256_256 vdd_d vss_d / DCAP4LVT
XXFILLER_256_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_257_256 vdd_d vss_d / DCAP4LVT
XXFILLER_257_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_258_256 vdd_d vss_d / DCAP4LVT
XXFILLER_258_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_259_256 vdd_d vss_d / DCAP4LVT
XXFILLER_259_2343 vdd_d vss_d / DCAP4LVT
XXFILLER_19_528 vdd_d vss_d / DCAP8LVT
XXFILLER_18_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_15_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_14_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_13_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_12_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_11_528 vdd_d vss_d / DCAP8LVT
XXFILLER_9_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_7_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_6_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_8_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_5_384 vdd_d vss_d / DCAP8LVT
XXFILLER_4_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_4_384 vdd_d vss_d / DCAP8LVT
XXFILLER_3_2340 vdd_d vss_d / DCAP8LVT
XXFILLER_2_2338 vdd_d vss_d / DCAP8LVT
XXFILLER_2_510 vdd_d vss_d / DCAP8LVT
XXFILLER_2_804 vdd_d vss_d / DCAP8LVT
XXFILLER_2_526 vdd_d vss_d / DCAP8LVT
XXFILLER_2_607 vdd_d vss_d / DCAP8LVT
XXFILLER_1_2335 vdd_d vss_d / DCAP8LVT
XXFILLER_1_816 vdd_d vss_d / DCAP8LVT
XXFILLER_2_690 vdd_d vss_d / DCAP8LVT
XXFILLER_16_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_20_1024 vdd_d vss_d / DCAP8LVT
XXFILLER_19_2339 vdd_d vss_d / DCAP8LVT
XXFILLER_0_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_20_1151 vdd_d vss_d / DCAP8LVT
XXFILLER_20_1604 vdd_d vss_d / DCAP8LVT
XXFILLER_20_1708 vdd_d vss_d / DCAP8LVT
XXFILLER_20_1742 vdd_d vss_d / DCAP8LVT
XXFILLER_20_2338 vdd_d vss_d / DCAP8LVT
XXFILLER_21_1142 vdd_d vss_d / DCAP8LVT
XXFILLER_21_1166 vdd_d vss_d / DCAP8LVT
XXFILLER_21_1216 vdd_d vss_d / DCAP8LVT
XXFILLER_21_1235 vdd_d vss_d / DCAP8LVT
XXFILLER_21_1597 vdd_d vss_d / DCAP8LVT
XXFILLER_22_1130 vdd_d vss_d / DCAP8LVT
XXFILLER_22_1148 vdd_d vss_d / DCAP8LVT
XXFILLER_22_1224 vdd_d vss_d / DCAP8LVT
XXFILLER_23_432 vdd_d vss_d / DCAP8LVT
XXFILLER_23_1037 vdd_d vss_d / DCAP8LVT
XXFILLER_23_1099 vdd_d vss_d / DCAP8LVT
XXFILLER_23_1111 vdd_d vss_d / DCAP8LVT
XXFILLER_23_1186 vdd_d vss_d / DCAP8LVT
XXFILLER_23_1218 vdd_d vss_d / DCAP8LVT
XXFILLER_23_1237 vdd_d vss_d / DCAP8LVT
XXFILLER_23_2337 vdd_d vss_d / DCAP8LVT
XXFILLER_24_1652 vdd_d vss_d / DCAP8LVT
XXFILLER_24_2341 vdd_d vss_d / DCAP8LVT
XXFILLER_25_512 vdd_d vss_d / DCAP8LVT
XXFILLER_25_1040 vdd_d vss_d / DCAP8LVT
XXFILLER_25_1109 vdd_d vss_d / DCAP8LVT
XXFILLER_25_1145 vdd_d vss_d / DCAP8LVT
XXFILLER_25_1160 vdd_d vss_d / DCAP8LVT
XXFILLER_25_1279 vdd_d vss_d / DCAP8LVT
XXFILLER_26_384 vdd_d vss_d / DCAP8LVT
XXFILLER_26_434 vdd_d vss_d / DCAP8LVT
XXFILLER_26_1035 vdd_d vss_d / DCAP8LVT
XXFILLER_26_1061 vdd_d vss_d / DCAP8LVT
XXFILLER_26_1217 vdd_d vss_d / DCAP8LVT
XXFILLER_26_1723 vdd_d vss_d / DCAP8LVT
XXFILLER_27_952 vdd_d vss_d / DCAP8LVT
XXFILLER_27_1024 vdd_d vss_d / DCAP8LVT
XXFILLER_27_1794 vdd_d vss_d / DCAP8LVT
XXFILLER_27_1825 vdd_d vss_d / DCAP8LVT
XXFILLER_27_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_28_432 vdd_d vss_d / DCAP8LVT
XXFILLER_28_585 vdd_d vss_d / DCAP8LVT
XXFILLER_28_894 vdd_d vss_d / DCAP8LVT
XXFILLER_28_1233 vdd_d vss_d / DCAP8LVT
XXFILLER_28_2337 vdd_d vss_d / DCAP8LVT
XXFILLER_29_432 vdd_d vss_d / DCAP8LVT
XXFILLER_29_1013 vdd_d vss_d / DCAP8LVT
XXFILLER_29_1172 vdd_d vss_d / DCAP8LVT
XXFILLER_29_1839 vdd_d vss_d / DCAP8LVT
XXFILLER_29_2335 vdd_d vss_d / DCAP8LVT
XXFILLER_30_416 vdd_d vss_d / DCAP8LVT
XXFILLER_30_1788 vdd_d vss_d / DCAP8LVT
XXFILLER_31_422 vdd_d vss_d / DCAP8LVT
XXFILLER_31_774 vdd_d vss_d / DCAP8LVT
XXFILLER_31_1864 vdd_d vss_d / DCAP8LVT
XXFILLER_31_2340 vdd_d vss_d / DCAP8LVT
XXFILLER_32_406 vdd_d vss_d / DCAP8LVT
XXFILLER_32_780 vdd_d vss_d / DCAP8LVT
XXFILLER_32_1094 vdd_d vss_d / DCAP8LVT
XXFILLER_32_1461 vdd_d vss_d / DCAP8LVT
XXFILLER_32_2342 vdd_d vss_d / DCAP8LVT
XXFILLER_33_457 vdd_d vss_d / DCAP8LVT
XXFILLER_33_1327 vdd_d vss_d / DCAP8LVT
XXFILLER_33_1407 vdd_d vss_d / DCAP8LVT
XXFILLER_33_2335 vdd_d vss_d / DCAP8LVT
XXFILLER_34_400 vdd_d vss_d / DCAP8LVT
XXFILLER_34_417 vdd_d vss_d / DCAP8LVT
XXFILLER_34_988 vdd_d vss_d / DCAP8LVT
XXFILLER_34_1083 vdd_d vss_d / DCAP8LVT
XXFILLER_34_1130 vdd_d vss_d / DCAP8LVT
XXFILLER_34_2335 vdd_d vss_d / DCAP8LVT
XXFILLER_35_499 vdd_d vss_d / DCAP8LVT
XXFILLER_35_572 vdd_d vss_d / DCAP8LVT
XXFILLER_35_1215 vdd_d vss_d / DCAP8LVT
XXFILLER_35_1291 vdd_d vss_d / DCAP8LVT
XXFILLER_35_1472 vdd_d vss_d / DCAP8LVT
XXFILLER_35_1542 vdd_d vss_d / DCAP8LVT
XXFILLER_36_400 vdd_d vss_d / DCAP8LVT
XXFILLER_36_850 vdd_d vss_d / DCAP8LVT
XXFILLER_36_1023 vdd_d vss_d / DCAP8LVT
XXFILLER_36_1068 vdd_d vss_d / DCAP8LVT
XXFILLER_36_1272 vdd_d vss_d / DCAP8LVT
XXFILLER_36_1396 vdd_d vss_d / DCAP8LVT
XXFILLER_36_1416 vdd_d vss_d / DCAP8LVT
XXFILLER_36_1451 vdd_d vss_d / DCAP8LVT
XXFILLER_36_1785 vdd_d vss_d / DCAP8LVT
XXFILLER_36_1872 vdd_d vss_d / DCAP8LVT
XXFILLER_36_2340 vdd_d vss_d / DCAP8LVT
XXFILLER_37_525 vdd_d vss_d / DCAP8LVT
XXFILLER_37_821 vdd_d vss_d / DCAP8LVT
XXFILLER_37_885 vdd_d vss_d / DCAP8LVT
XXFILLER_37_1675 vdd_d vss_d / DCAP8LVT
XXFILLER_37_1820 vdd_d vss_d / DCAP8LVT
XXFILLER_37_1904 vdd_d vss_d / DCAP8LVT
XXFILLER_38_416 vdd_d vss_d / DCAP8LVT
XXFILLER_38_447 vdd_d vss_d / DCAP8LVT
XXFILLER_38_756 vdd_d vss_d / DCAP8LVT
XXFILLER_38_800 vdd_d vss_d / DCAP8LVT
XXFILLER_38_1067 vdd_d vss_d / DCAP8LVT
XXFILLER_38_1089 vdd_d vss_d / DCAP8LVT
XXFILLER_38_1189 vdd_d vss_d / DCAP8LVT
XXFILLER_38_1345 vdd_d vss_d / DCAP8LVT
XXFILLER_38_1443 vdd_d vss_d / DCAP8LVT
XXFILLER_38_1546 vdd_d vss_d / DCAP8LVT
XXFILLER_38_1732 vdd_d vss_d / DCAP8LVT
XXFILLER_38_1796 vdd_d vss_d / DCAP8LVT
XXFILLER_38_1837 vdd_d vss_d / DCAP8LVT
XXFILLER_38_2338 vdd_d vss_d / DCAP8LVT
XXFILLER_39_506 vdd_d vss_d / DCAP8LVT
XXFILLER_39_744 vdd_d vss_d / DCAP8LVT
XXFILLER_39_941 vdd_d vss_d / DCAP8LVT
XXFILLER_39_1235 vdd_d vss_d / DCAP8LVT
XXFILLER_39_1276 vdd_d vss_d / DCAP8LVT
XXFILLER_39_1370 vdd_d vss_d / DCAP8LVT
XXFILLER_39_1419 vdd_d vss_d / DCAP8LVT
XXFILLER_39_1470 vdd_d vss_d / DCAP8LVT
XXFILLER_39_1575 vdd_d vss_d / DCAP8LVT
XXFILLER_39_1816 vdd_d vss_d / DCAP8LVT
XXFILLER_40_425 vdd_d vss_d / DCAP8LVT
XXFILLER_40_611 vdd_d vss_d / DCAP8LVT
XXFILLER_40_721 vdd_d vss_d / DCAP8LVT
XXFILLER_40_778 vdd_d vss_d / DCAP8LVT
XXFILLER_40_895 vdd_d vss_d / DCAP8LVT
XXFILLER_40_951 vdd_d vss_d / DCAP8LVT
XXFILLER_40_966 vdd_d vss_d / DCAP8LVT
XXFILLER_40_1374 vdd_d vss_d / DCAP8LVT
XXFILLER_41_384 vdd_d vss_d / DCAP8LVT
XXFILLER_41_430 vdd_d vss_d / DCAP8LVT
XXFILLER_41_816 vdd_d vss_d / DCAP8LVT
XXFILLER_41_838 vdd_d vss_d / DCAP8LVT
XXFILLER_41_945 vdd_d vss_d / DCAP8LVT
XXFILLER_41_1036 vdd_d vss_d / DCAP8LVT
XXFILLER_41_1136 vdd_d vss_d / DCAP8LVT
XXFILLER_41_1237 vdd_d vss_d / DCAP8LVT
XXFILLER_41_1492 vdd_d vss_d / DCAP8LVT
XXFILLER_41_1586 vdd_d vss_d / DCAP8LVT
XXFILLER_41_1859 vdd_d vss_d / DCAP8LVT
XXFILLER_41_2339 vdd_d vss_d / DCAP8LVT
XXFILLER_42_384 vdd_d vss_d / DCAP8LVT
XXFILLER_42_703 vdd_d vss_d / DCAP8LVT
XXFILLER_42_747 vdd_d vss_d / DCAP8LVT
XXFILLER_42_813 vdd_d vss_d / DCAP8LVT
XXFILLER_42_852 vdd_d vss_d / DCAP8LVT
XXFILLER_42_890 vdd_d vss_d / DCAP8LVT
XXFILLER_42_912 vdd_d vss_d / DCAP8LVT
XXFILLER_42_975 vdd_d vss_d / DCAP8LVT
XXFILLER_42_1111 vdd_d vss_d / DCAP8LVT
XXFILLER_42_1209 vdd_d vss_d / DCAP8LVT
XXFILLER_42_1319 vdd_d vss_d / DCAP8LVT
XXFILLER_42_1415 vdd_d vss_d / DCAP8LVT
XXFILLER_42_1503 vdd_d vss_d / DCAP8LVT
XXFILLER_42_1533 vdd_d vss_d / DCAP8LVT
XXFILLER_42_1553 vdd_d vss_d / DCAP8LVT
XXFILLER_42_1655 vdd_d vss_d / DCAP8LVT
XXFILLER_42_1906 vdd_d vss_d / DCAP8LVT
XXFILLER_42_1994 vdd_d vss_d / DCAP8LVT
XXFILLER_43_493 vdd_d vss_d / DCAP8LVT
XXFILLER_43_786 vdd_d vss_d / DCAP8LVT
XXFILLER_43_1103 vdd_d vss_d / DCAP8LVT
XXFILLER_43_1357 vdd_d vss_d / DCAP8LVT
XXFILLER_43_1639 vdd_d vss_d / DCAP8LVT
XXFILLER_43_1793 vdd_d vss_d / DCAP8LVT
XXFILLER_43_1829 vdd_d vss_d / DCAP8LVT
XXFILLER_43_1878 vdd_d vss_d / DCAP8LVT
XXFILLER_43_1942 vdd_d vss_d / DCAP8LVT
XXFILLER_43_2338 vdd_d vss_d / DCAP8LVT
XXFILLER_44_375 vdd_d vss_d / DCAP8LVT
XXFILLER_44_436 vdd_d vss_d / DCAP8LVT
XXFILLER_44_454 vdd_d vss_d / DCAP8LVT
XXFILLER_44_802 vdd_d vss_d / DCAP8LVT
XXFILLER_44_890 vdd_d vss_d / DCAP8LVT
XXFILLER_44_904 vdd_d vss_d / DCAP8LVT
XXFILLER_44_1143 vdd_d vss_d / DCAP8LVT
XXFILLER_44_1211 vdd_d vss_d / DCAP8LVT
XXFILLER_44_1361 vdd_d vss_d / DCAP8LVT
XXFILLER_44_1502 vdd_d vss_d / DCAP8LVT
XXFILLER_44_1525 vdd_d vss_d / DCAP8LVT
XXFILLER_44_1561 vdd_d vss_d / DCAP8LVT
XXFILLER_44_1581 vdd_d vss_d / DCAP8LVT
XXFILLER_44_1601 vdd_d vss_d / DCAP8LVT
XXFILLER_44_1624 vdd_d vss_d / DCAP8LVT
XXFILLER_44_1716 vdd_d vss_d / DCAP8LVT
XXFILLER_44_1910 vdd_d vss_d / DCAP8LVT
XXFILLER_45_720 vdd_d vss_d / DCAP8LVT
XXFILLER_45_924 vdd_d vss_d / DCAP8LVT
XXFILLER_45_2339 vdd_d vss_d / DCAP8LVT
XXFILLER_46_896 vdd_d vss_d / DCAP8LVT
XXFILLER_46_1680 vdd_d vss_d / DCAP8LVT
XXFILLER_46_2335 vdd_d vss_d / DCAP8LVT
XXFILLER_47_656 vdd_d vss_d / DCAP8LVT
XXFILLER_48_80 vdd_d vss_d / DCAP8LVT
XXFILLER_48_2253 vdd_d vss_d / DCAP8LVT
XXFILLER_48_2335 vdd_d vss_d / DCAP8LVT
XXFILLER_49_400 vdd_d vss_d / DCAP8LVT
XXFILLER_49_1479 vdd_d vss_d / DCAP8LVT
XXFILLER_49_2337 vdd_d vss_d / DCAP8LVT
XXFILLER_50_384 vdd_d vss_d / DCAP8LVT
XXFILLER_50_402 vdd_d vss_d / DCAP8LVT
XXFILLER_50_811 vdd_d vss_d / DCAP8LVT
XXFILLER_50_1729 vdd_d vss_d / DCAP8LVT
XXFILLER_51_1248 vdd_d vss_d / DCAP8LVT
XXFILLER_52_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_53_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_54_893 vdd_d vss_d / DCAP8LVT
XXFILLER_55_416 vdd_d vss_d / DCAP8LVT
XXFILLER_55_1936 vdd_d vss_d / DCAP8LVT
XXFILLER_57_1753 vdd_d vss_d / DCAP8LVT
XXFILLER_65_747 vdd_d vss_d / DCAP8LVT
XXFILLER_66_715 vdd_d vss_d / DCAP8LVT
XXFILLER_68_1253 vdd_d vss_d / DCAP8LVT
XXFILLER_72_1103 vdd_d vss_d / DCAP8LVT
XXFILLER_72_1248 vdd_d vss_d / DCAP8LVT
XXFILLER_73_240 vdd_d vss_d / DCAP8LVT
XXFILLER_74_1119 vdd_d vss_d / DCAP8LVT
XXFILLER_74_1249 vdd_d vss_d / DCAP8LVT
XXFILLER_76_240 vdd_d vss_d / DCAP8LVT
XXFILLER_77_1199 vdd_d vss_d / DCAP8LVT
XXFILLER_82_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_83_1231 vdd_d vss_d / DCAP8LVT
XXFILLER_83_1250 vdd_d vss_d / DCAP8LVT
XXFILLER_85_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_92_1215 vdd_d vss_d / DCAP8LVT
XXFILLER_93_1731 vdd_d vss_d / DCAP8LVT
XXFILLER_95_400 vdd_d vss_d / DCAP8LVT
XXFILLER_95_439 vdd_d vss_d / DCAP8LVT
XXFILLER_95_949 vdd_d vss_d / DCAP8LVT
XXFILLER_95_1404 vdd_d vss_d / DCAP8LVT
XXFILLER_96_352 vdd_d vss_d / DCAP8LVT
XXFILLER_96_401 vdd_d vss_d / DCAP8LVT
XXFILLER_96_1371 vdd_d vss_d / DCAP8LVT
XXFILLER_96_2340 vdd_d vss_d / DCAP8LVT
XXFILLER_97_336 vdd_d vss_d / DCAP8LVT
XXFILLER_97_449 vdd_d vss_d / DCAP8LVT
XXFILLER_97_2342 vdd_d vss_d / DCAP8LVT
XXFILLER_98_1609 vdd_d vss_d / DCAP8LVT
XXFILLER_98_2340 vdd_d vss_d / DCAP8LVT
XXFILLER_99_1406 vdd_d vss_d / DCAP8LVT
XXFILLER_99_1906 vdd_d vss_d / DCAP8LVT
XXFILLER_100_1168 vdd_d vss_d / DCAP8LVT
XXFILLER_101_1949 vdd_d vss_d / DCAP8LVT
XXFILLER_101_2340 vdd_d vss_d / DCAP8LVT
XXFILLER_102_1024 vdd_d vss_d / DCAP8LVT
XXFILLER_102_2340 vdd_d vss_d / DCAP8LVT
XXFILLER_103_1900 vdd_d vss_d / DCAP8LVT
XXFILLER_104_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_105_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_106_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_107_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_108_1406 vdd_d vss_d / DCAP8LVT
XXFILLER_108_2339 vdd_d vss_d / DCAP8LVT
XXFILLER_109_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_110_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_111_1857 vdd_d vss_d / DCAP8LVT
XXFILLER_131_240 vdd_d vss_d / DCAP8LVT
XXFILLER_131_2339 vdd_d vss_d / DCAP8LVT
XXFILLER_136_748 vdd_d vss_d / DCAP8LVT
XXFILLER_136_1749 vdd_d vss_d / DCAP8LVT
XXFILLER_140_1167 vdd_d vss_d / DCAP8LVT
XXFILLER_150_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_151_432 vdd_d vss_d / DCAP8LVT
XXFILLER_151_936 vdd_d vss_d / DCAP8LVT
XXFILLER_151_954 vdd_d vss_d / DCAP8LVT
XXFILLER_151_1407 vdd_d vss_d / DCAP8LVT
XXFILLER_152_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_153_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_154_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_155_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_156_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_157_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_158_2338 vdd_d vss_d / DCAP8LVT
XXFILLER_159_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_160_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_161_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_162_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_163_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_164_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_165_1856 vdd_d vss_d / DCAP8LVT
XXFILLER_165_2337 vdd_d vss_d / DCAP8LVT
XXFILLER_166_1406 vdd_d vss_d / DCAP8LVT
XXFILLER_166_1874 vdd_d vss_d / DCAP8LVT
XXFILLER_180_1167 vdd_d vss_d / DCAP8LVT
XXFILLER_181_1144 vdd_d vss_d / DCAP8LVT
XXFILLER_181_1245 vdd_d vss_d / DCAP8LVT
XXFILLER_182_1230 vdd_d vss_d / DCAP8LVT
XXFILLER_183_1240 vdd_d vss_d / DCAP8LVT
XXFILLER_206_1420 vdd_d vss_d / DCAP8LVT
XXFILLER_206_2340 vdd_d vss_d / DCAP8LVT
XXFILLER_207_928 vdd_d vss_d / DCAP8LVT
XXFILLER_207_2342 vdd_d vss_d / DCAP8LVT
XXFILLER_208_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_209_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_210_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_211_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_212_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_213_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_214_688 vdd_d vss_d / DCAP8LVT
XXFILLER_214_2337 vdd_d vss_d / DCAP8LVT
XXFILLER_215_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_216_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_217_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_218_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_219_896 vdd_d vss_d / DCAP8LVT
XXFILLER_219_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_220_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_221_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_222_2336 vdd_d vss_d / DCAP8LVT
XXFILLER_19_512 vdd_d vss_d / DCAP16LVT
XXFILLER_11_2334 vdd_d vss_d / DCAP16LVT
XXFILLER_11_512 vdd_d vss_d / DCAP16LVT
XXFILLER_10_800 vdd_d vss_d / DCAP16LVT
XXFILLER_5_2331 vdd_d vss_d / DCAP16LVT
XXFILLER_3_395 vdd_d vss_d / DCAP16LVT
XXFILLER_2_761 vdd_d vss_d / DCAP16LVT
XXFILLER_2_494 vdd_d vss_d / DCAP16LVT
XXFILLER_2_788 vdd_d vss_d / DCAP16LVT
XXFILLER_2_733 vdd_d vss_d / DCAP16LVT
XXFILLER_1_800 vdd_d vss_d / DCAP16LVT
XXFILLER_20_1135 vdd_d vss_d / DCAP16LVT
XXFILLER_19_2323 vdd_d vss_d / DCAP16LVT
XXFILLER_20_1692 vdd_d vss_d / DCAP16LVT
XXFILLER_20_1726 vdd_d vss_d / DCAP16LVT
XXFILLER_21_448 vdd_d vss_d / DCAP16LVT
XXFILLER_21_1581 vdd_d vss_d / DCAP16LVT
XXFILLER_22_1310 vdd_d vss_d / DCAP16LVT
XXFILLER_22_2327 vdd_d vss_d / DCAP16LVT
XXFILLER_23_416 vdd_d vss_d / DCAP16LVT
XXFILLER_23_1083 vdd_d vss_d / DCAP16LVT
XXFILLER_23_1170 vdd_d vss_d / DCAP16LVT
XXFILLER_23_1202 vdd_d vss_d / DCAP16LVT
XXFILLER_23_1748 vdd_d vss_d / DCAP16LVT
XXFILLER_23_2321 vdd_d vss_d / DCAP16LVT
XXFILLER_24_384 vdd_d vss_d / DCAP16LVT
XXFILLER_24_1210 vdd_d vss_d / DCAP16LVT
XXFILLER_25_1129 vdd_d vss_d / DCAP16LVT
XXFILLER_25_1209 vdd_d vss_d / DCAP16LVT
XXFILLER_26_1406 vdd_d vss_d / DCAP16LVT
XXFILLER_27_384 vdd_d vss_d / DCAP16LVT
XXFILLER_27_479 vdd_d vss_d / DCAP16LVT
XXFILLER_27_1008 vdd_d vss_d / DCAP16LVT
XXFILLER_27_1778 vdd_d vss_d / DCAP16LVT
XXFILLER_27_1809 vdd_d vss_d / DCAP16LVT
XXFILLER_27_2320 vdd_d vss_d / DCAP16LVT
XXFILLER_28_461 vdd_d vss_d / DCAP16LVT
XXFILLER_28_496 vdd_d vss_d / DCAP16LVT
XXFILLER_28_1217 vdd_d vss_d / DCAP16LVT
XXFILLER_29_416 vdd_d vss_d / DCAP16LVT
XXFILLER_29_997 vdd_d vss_d / DCAP16LVT
XXFILLER_29_1156 vdd_d vss_d / DCAP16LVT
XXFILLER_29_1317 vdd_d vss_d / DCAP16LVT
XXFILLER_29_1823 vdd_d vss_d / DCAP16LVT
XXFILLER_30_978 vdd_d vss_d / DCAP16LVT
XXFILLER_30_1772 vdd_d vss_d / DCAP16LVT
XXFILLER_31_465 vdd_d vss_d / DCAP16LVT
XXFILLER_31_1848 vdd_d vss_d / DCAP16LVT
XXFILLER_32_390 vdd_d vss_d / DCAP16LVT
XXFILLER_32_966 vdd_d vss_d / DCAP16LVT
XXFILLER_32_1403 vdd_d vss_d / DCAP16LVT
XXFILLER_32_1837 vdd_d vss_d / DCAP16LVT
XXFILLER_33_1127 vdd_d vss_d / DCAP16LVT
XXFILLER_33_1783 vdd_d vss_d / DCAP16LVT
XXFILLER_33_2319 vdd_d vss_d / DCAP16LVT
XXFILLER_34_384 vdd_d vss_d / DCAP16LVT
XXFILLER_34_1067 vdd_d vss_d / DCAP16LVT
XXFILLER_34_1401 vdd_d vss_d / DCAP16LVT
XXFILLER_34_1490 vdd_d vss_d / DCAP16LVT
XXFILLER_35_1199 vdd_d vss_d / DCAP16LVT
XXFILLER_35_1405 vdd_d vss_d / DCAP16LVT
XXFILLER_35_1526 vdd_d vss_d / DCAP16LVT
XXFILLER_35_2331 vdd_d vss_d / DCAP16LVT
XXFILLER_36_384 vdd_d vss_d / DCAP16LVT
XXFILLER_36_739 vdd_d vss_d / DCAP16LVT
XXFILLER_36_793 vdd_d vss_d / DCAP16LVT
XXFILLER_36_1244 vdd_d vss_d / DCAP16LVT
XXFILLER_36_1435 vdd_d vss_d / DCAP16LVT
XXFILLER_37_461 vdd_d vss_d / DCAP16LVT
XXFILLER_37_805 vdd_d vss_d / DCAP16LVT
XXFILLER_37_869 vdd_d vss_d / DCAP16LVT
XXFILLER_37_1133 vdd_d vss_d / DCAP16LVT
XXFILLER_37_1187 vdd_d vss_d / DCAP16LVT
XXFILLER_37_1309 vdd_d vss_d / DCAP16LVT
XXFILLER_38_431 vdd_d vss_d / DCAP16LVT
XXFILLER_38_621 vdd_d vss_d / DCAP16LVT
XXFILLER_38_740 vdd_d vss_d / DCAP16LVT
XXFILLER_38_849 vdd_d vss_d / DCAP16LVT
XXFILLER_38_1007 vdd_d vss_d / DCAP16LVT
XXFILLER_38_1427 vdd_d vss_d / DCAP16LVT
XXFILLER_38_1491 vdd_d vss_d / DCAP16LVT
XXFILLER_38_1780 vdd_d vss_d / DCAP16LVT
XXFILLER_38_1821 vdd_d vss_d / DCAP16LVT
XXFILLER_38_1918 vdd_d vss_d / DCAP16LVT
XXFILLER_38_2322 vdd_d vss_d / DCAP16LVT
XXFILLER_39_826 vdd_d vss_d / DCAP16LVT
XXFILLER_39_989 vdd_d vss_d / DCAP16LVT
XXFILLER_39_1354 vdd_d vss_d / DCAP16LVT
XXFILLER_39_1517 vdd_d vss_d / DCAP16LVT
XXFILLER_39_2328 vdd_d vss_d / DCAP16LVT
XXFILLER_40_558 vdd_d vss_d / DCAP16LVT
XXFILLER_40_879 vdd_d vss_d / DCAP16LVT
XXFILLER_40_926 vdd_d vss_d / DCAP16LVT
XXFILLER_40_1038 vdd_d vss_d / DCAP16LVT
XXFILLER_40_1096 vdd_d vss_d / DCAP16LVT
XXFILLER_40_1153 vdd_d vss_d / DCAP16LVT
XXFILLER_40_1639 vdd_d vss_d / DCAP16LVT
XXFILLER_40_1755 vdd_d vss_d / DCAP16LVT
XXFILLER_41_800 vdd_d vss_d / DCAP16LVT
XXFILLER_41_862 vdd_d vss_d / DCAP16LVT
XXFILLER_41_929 vdd_d vss_d / DCAP16LVT
XXFILLER_41_1120 vdd_d vss_d / DCAP16LVT
XXFILLER_41_1156 vdd_d vss_d / DCAP16LVT
XXFILLER_41_1570 vdd_d vss_d / DCAP16LVT
XXFILLER_41_1686 vdd_d vss_d / DCAP16LVT
XXFILLER_42_550 vdd_d vss_d / DCAP16LVT
XXFILLER_42_1081 vdd_d vss_d / DCAP16LVT
XXFILLER_42_1338 vdd_d vss_d / DCAP16LVT
XXFILLER_42_1487 vdd_d vss_d / DCAP16LVT
XXFILLER_42_1639 vdd_d vss_d / DCAP16LVT
XXFILLER_42_1797 vdd_d vss_d / DCAP16LVT
XXFILLER_42_1978 vdd_d vss_d / DCAP16LVT
XXFILLER_42_2328 vdd_d vss_d / DCAP16LVT
XXFILLER_43_756 vdd_d vss_d / DCAP16LVT
XXFILLER_43_866 vdd_d vss_d / DCAP16LVT
XXFILLER_43_934 vdd_d vss_d / DCAP16LVT
XXFILLER_43_1295 vdd_d vss_d / DCAP16LVT
XXFILLER_43_1475 vdd_d vss_d / DCAP16LVT
XXFILLER_43_1521 vdd_d vss_d / DCAP16LVT
XXFILLER_43_1777 vdd_d vss_d / DCAP16LVT
XXFILLER_43_1813 vdd_d vss_d / DCAP16LVT
XXFILLER_43_1926 vdd_d vss_d / DCAP16LVT
XXFILLER_44_352 vdd_d vss_d / DCAP16LVT
XXFILLER_44_758 vdd_d vss_d / DCAP16LVT
XXFILLER_44_874 vdd_d vss_d / DCAP16LVT
XXFILLER_44_986 vdd_d vss_d / DCAP16LVT
XXFILLER_44_1067 vdd_d vss_d / DCAP16LVT
XXFILLER_44_1168 vdd_d vss_d / DCAP16LVT
XXFILLER_44_1345 vdd_d vss_d / DCAP16LVT
XXFILLER_44_1382 vdd_d vss_d / DCAP16LVT
XXFILLER_44_1407 vdd_d vss_d / DCAP16LVT
XXFILLER_44_1461 vdd_d vss_d / DCAP16LVT
XXFILLER_44_1639 vdd_d vss_d / DCAP16LVT
XXFILLER_44_1817 vdd_d vss_d / DCAP16LVT
XXFILLER_44_1846 vdd_d vss_d / DCAP16LVT
XXFILLER_44_1871 vdd_d vss_d / DCAP16LVT
XXFILLER_44_2330 vdd_d vss_d / DCAP16LVT
XXFILLER_45_704 vdd_d vss_d / DCAP16LVT
XXFILLER_45_1573 vdd_d vss_d / DCAP16LVT
XXFILLER_45_1878 vdd_d vss_d / DCAP16LVT
XXFILLER_45_2323 vdd_d vss_d / DCAP16LVT
XXFILLER_46_1937 vdd_d vss_d / DCAP16LVT
XXFILLER_47_640 vdd_d vss_d / DCAP16LVT
XXFILLER_48_64 vdd_d vss_d / DCAP16LVT
XXFILLER_48_2237 vdd_d vss_d / DCAP16LVT
XXFILLER_49_384 vdd_d vss_d / DCAP16LVT
XXFILLER_49_2321 vdd_d vss_d / DCAP16LVT
XXFILLER_50_795 vdd_d vss_d / DCAP16LVT
XXFILLER_50_1469 vdd_d vss_d / DCAP16LVT
XXFILLER_50_1713 vdd_d vss_d / DCAP16LVT
XXFILLER_50_1898 vdd_d vss_d / DCAP16LVT
XXFILLER_50_2334 vdd_d vss_d / DCAP16LVT
XXFILLER_53_1184 vdd_d vss_d / DCAP16LVT
XXFILLER_53_2320 vdd_d vss_d / DCAP16LVT
XXFILLER_54_800 vdd_d vss_d / DCAP16LVT
XXFILLER_54_1927 vdd_d vss_d / DCAP16LVT
XXFILLER_55_2330 vdd_d vss_d / DCAP16LVT
XXFILLER_56_747 vdd_d vss_d / DCAP16LVT
XXFILLER_56_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_56_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_57_747 vdd_d vss_d / DCAP16LVT
XXFILLER_57_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_57_1651 vdd_d vss_d / DCAP16LVT
XXFILLER_57_1737 vdd_d vss_d / DCAP16LVT
XXFILLER_58_747 vdd_d vss_d / DCAP16LVT
XXFILLER_58_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_58_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_59_747 vdd_d vss_d / DCAP16LVT
XXFILLER_59_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_59_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_60_747 vdd_d vss_d / DCAP16LVT
XXFILLER_60_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_60_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_61_747 vdd_d vss_d / DCAP16LVT
XXFILLER_61_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_61_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_62_747 vdd_d vss_d / DCAP16LVT
XXFILLER_62_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_62_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_63_747 vdd_d vss_d / DCAP16LVT
XXFILLER_63_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_63_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_64_747 vdd_d vss_d / DCAP16LVT
XXFILLER_64_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_64_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_65_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_65_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_66_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_66_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_67_747 vdd_d vss_d / DCAP16LVT
XXFILLER_67_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_67_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_68_747 vdd_d vss_d / DCAP16LVT
XXFILLER_68_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_69_224 vdd_d vss_d / DCAP16LVT
XXFILLER_69_747 vdd_d vss_d / DCAP16LVT
XXFILLER_69_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_69_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_69_2327 vdd_d vss_d / DCAP16LVT
XXFILLER_70_747 vdd_d vss_d / DCAP16LVT
XXFILLER_70_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_70_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_71_747 vdd_d vss_d / DCAP16LVT
XXFILLER_71_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_71_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_72_747 vdd_d vss_d / DCAP16LVT
XXFILLER_72_1087 vdd_d vss_d / DCAP16LVT
XXFILLER_72_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_73_224 vdd_d vss_d / DCAP16LVT
XXFILLER_73_747 vdd_d vss_d / DCAP16LVT
XXFILLER_73_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_73_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_74_747 vdd_d vss_d / DCAP16LVT
XXFILLER_74_1233 vdd_d vss_d / DCAP16LVT
XXFILLER_74_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_75_747 vdd_d vss_d / DCAP16LVT
XXFILLER_75_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_76_224 vdd_d vss_d / DCAP16LVT
XXFILLER_76_747 vdd_d vss_d / DCAP16LVT
XXFILLER_76_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_76_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_77_747 vdd_d vss_d / DCAP16LVT
XXFILLER_77_1183 vdd_d vss_d / DCAP16LVT
XXFILLER_77_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_77_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_78_747 vdd_d vss_d / DCAP16LVT
XXFILLER_78_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_78_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_79_747 vdd_d vss_d / DCAP16LVT
XXFILLER_79_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_79_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_80_747 vdd_d vss_d / DCAP16LVT
XXFILLER_80_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_80_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_81_747 vdd_d vss_d / DCAP16LVT
XXFILLER_81_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_81_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_82_747 vdd_d vss_d / DCAP16LVT
XXFILLER_82_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_82_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_82_2320 vdd_d vss_d / DCAP16LVT
XXFILLER_83_747 vdd_d vss_d / DCAP16LVT
XXFILLER_83_1215 vdd_d vss_d / DCAP16LVT
XXFILLER_83_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_84_747 vdd_d vss_d / DCAP16LVT
XXFILLER_84_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_84_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_85_747 vdd_d vss_d / DCAP16LVT
XXFILLER_85_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_85_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_85_2320 vdd_d vss_d / DCAP16LVT
XXFILLER_86_747 vdd_d vss_d / DCAP16LVT
XXFILLER_86_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_86_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_87_747 vdd_d vss_d / DCAP16LVT
XXFILLER_87_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_87_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_88_747 vdd_d vss_d / DCAP16LVT
XXFILLER_88_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_88_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_89_747 vdd_d vss_d / DCAP16LVT
XXFILLER_89_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_89_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_90_747 vdd_d vss_d / DCAP16LVT
XXFILLER_90_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_90_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_91_747 vdd_d vss_d / DCAP16LVT
XXFILLER_91_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_91_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_92_747 vdd_d vss_d / DCAP16LVT
XXFILLER_92_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_93_747 vdd_d vss_d / DCAP16LVT
XXFILLER_93_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_93_1715 vdd_d vss_d / DCAP16LVT
XXFILLER_94_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_94_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_95_384 vdd_d vss_d / DCAP16LVT
XXFILLER_95_423 vdd_d vss_d / DCAP16LVT
XXFILLER_95_923 vdd_d vss_d / DCAP16LVT
XXFILLER_95_1867 vdd_d vss_d / DCAP16LVT
XXFILLER_96_1355 vdd_d vss_d / DCAP16LVT
XXFILLER_96_2324 vdd_d vss_d / DCAP16LVT
XXFILLER_97_320 vdd_d vss_d / DCAP16LVT
XXFILLER_97_1430 vdd_d vss_d / DCAP16LVT
XXFILLER_97_2326 vdd_d vss_d / DCAP16LVT
XXFILLER_98_1788 vdd_d vss_d / DCAP16LVT
XXFILLER_98_2324 vdd_d vss_d / DCAP16LVT
XXFILLER_99_960 vdd_d vss_d / DCAP16LVT
XXFILLER_100_1152 vdd_d vss_d / DCAP16LVT
XXFILLER_100_2328 vdd_d vss_d / DCAP16LVT
XXFILLER_101_2324 vdd_d vss_d / DCAP16LVT
XXFILLER_102_1008 vdd_d vss_d / DCAP16LVT
XXFILLER_102_1294 vdd_d vss_d / DCAP16LVT
XXFILLER_103_1600 vdd_d vss_d / DCAP16LVT
XXFILLER_103_1884 vdd_d vss_d / DCAP16LVT
XXFILLER_103_2332 vdd_d vss_d / DCAP16LVT
XXFILLER_108_896 vdd_d vss_d / DCAP16LVT
XXFILLER_108_1390 vdd_d vss_d / DCAP16LVT
XXFILLER_111_1841 vdd_d vss_d / DCAP16LVT
XXFILLER_112_747 vdd_d vss_d / DCAP16LVT
XXFILLER_112_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_112_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_113_747 vdd_d vss_d / DCAP16LVT
XXFILLER_113_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_113_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_114_747 vdd_d vss_d / DCAP16LVT
XXFILLER_114_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_114_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_115_747 vdd_d vss_d / DCAP16LVT
XXFILLER_115_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_115_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_116_747 vdd_d vss_d / DCAP16LVT
XXFILLER_116_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_116_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_117_747 vdd_d vss_d / DCAP16LVT
XXFILLER_117_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_117_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_118_747 vdd_d vss_d / DCAP16LVT
XXFILLER_118_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_118_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_119_747 vdd_d vss_d / DCAP16LVT
XXFILLER_119_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_119_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_120_747 vdd_d vss_d / DCAP16LVT
XXFILLER_120_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_120_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_121_747 vdd_d vss_d / DCAP16LVT
XXFILLER_121_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_121_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_122_747 vdd_d vss_d / DCAP16LVT
XXFILLER_122_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_122_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_123_747 vdd_d vss_d / DCAP16LVT
XXFILLER_123_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_123_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_124_747 vdd_d vss_d / DCAP16LVT
XXFILLER_124_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_124_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_125_747 vdd_d vss_d / DCAP16LVT
XXFILLER_125_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_125_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_126_747 vdd_d vss_d / DCAP16LVT
XXFILLER_126_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_126_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_127_747 vdd_d vss_d / DCAP16LVT
XXFILLER_127_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_128_747 vdd_d vss_d / DCAP16LVT
XXFILLER_128_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_128_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_129_747 vdd_d vss_d / DCAP16LVT
XXFILLER_129_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_129_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_130_747 vdd_d vss_d / DCAP16LVT
XXFILLER_130_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_130_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_131_224 vdd_d vss_d / DCAP16LVT
XXFILLER_131_747 vdd_d vss_d / DCAP16LVT
XXFILLER_131_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_131_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_131_2323 vdd_d vss_d / DCAP16LVT
XXFILLER_132_747 vdd_d vss_d / DCAP16LVT
XXFILLER_132_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_132_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_133_747 vdd_d vss_d / DCAP16LVT
XXFILLER_133_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_133_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_134_747 vdd_d vss_d / DCAP16LVT
XXFILLER_134_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_134_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_135_747 vdd_d vss_d / DCAP16LVT
XXFILLER_135_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_135_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_136_715 vdd_d vss_d / DCAP16LVT
XXFILLER_136_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_136_1733 vdd_d vss_d / DCAP16LVT
XXFILLER_137_747 vdd_d vss_d / DCAP16LVT
XXFILLER_137_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_137_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_138_747 vdd_d vss_d / DCAP16LVT
XXFILLER_138_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_138_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_139_747 vdd_d vss_d / DCAP16LVT
XXFILLER_139_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_139_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_140_747 vdd_d vss_d / DCAP16LVT
XXFILLER_140_1151 vdd_d vss_d / DCAP16LVT
XXFILLER_140_1240 vdd_d vss_d / DCAP16LVT
XXFILLER_140_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_141_747 vdd_d vss_d / DCAP16LVT
XXFILLER_141_1246 vdd_d vss_d / DCAP16LVT
XXFILLER_141_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_142_747 vdd_d vss_d / DCAP16LVT
XXFILLER_142_1151 vdd_d vss_d / DCAP16LVT
XXFILLER_142_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_143_747 vdd_d vss_d / DCAP16LVT
XXFILLER_143_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_143_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_144_747 vdd_d vss_d / DCAP16LVT
XXFILLER_144_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_144_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_145_747 vdd_d vss_d / DCAP16LVT
XXFILLER_145_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_145_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_146_747 vdd_d vss_d / DCAP16LVT
XXFILLER_146_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_146_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_147_747 vdd_d vss_d / DCAP16LVT
XXFILLER_147_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_147_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_148_747 vdd_d vss_d / DCAP16LVT
XXFILLER_148_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_148_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_149_747 vdd_d vss_d / DCAP16LVT
XXFILLER_149_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_149_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_150_416 vdd_d vss_d / DCAP16LVT
XXFILLER_151_416 vdd_d vss_d / DCAP16LVT
XXFILLER_151_1391 vdd_d vss_d / DCAP16LVT
XXFILLER_158_672 vdd_d vss_d / DCAP16LVT
XXFILLER_166_896 vdd_d vss_d / DCAP16LVT
XXFILLER_166_1390 vdd_d vss_d / DCAP16LVT
XXFILLER_167_747 vdd_d vss_d / DCAP16LVT
XXFILLER_167_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_167_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_168_747 vdd_d vss_d / DCAP16LVT
XXFILLER_168_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_168_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_169_747 vdd_d vss_d / DCAP16LVT
XXFILLER_169_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_169_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_170_747 vdd_d vss_d / DCAP16LVT
XXFILLER_170_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_170_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_171_747 vdd_d vss_d / DCAP16LVT
XXFILLER_171_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_171_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_172_747 vdd_d vss_d / DCAP16LVT
XXFILLER_172_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_172_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_173_747 vdd_d vss_d / DCAP16LVT
XXFILLER_173_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_173_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_174_747 vdd_d vss_d / DCAP16LVT
XXFILLER_174_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_174_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_175_747 vdd_d vss_d / DCAP16LVT
XXFILLER_175_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_175_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_176_747 vdd_d vss_d / DCAP16LVT
XXFILLER_176_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_176_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_177_747 vdd_d vss_d / DCAP16LVT
XXFILLER_177_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_177_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_178_747 vdd_d vss_d / DCAP16LVT
XXFILLER_178_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_178_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_179_747 vdd_d vss_d / DCAP16LVT
XXFILLER_179_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_179_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_180_747 vdd_d vss_d / DCAP16LVT
XXFILLER_180_1151 vdd_d vss_d / DCAP16LVT
XXFILLER_180_1240 vdd_d vss_d / DCAP16LVT
XXFILLER_180_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_181_747 vdd_d vss_d / DCAP16LVT
XXFILLER_181_1128 vdd_d vss_d / DCAP16LVT
XXFILLER_181_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_182_747 vdd_d vss_d / DCAP16LVT
XXFILLER_182_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_183_747 vdd_d vss_d / DCAP16LVT
XXFILLER_183_1224 vdd_d vss_d / DCAP16LVT
XXFILLER_183_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_184_747 vdd_d vss_d / DCAP16LVT
XXFILLER_184_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_184_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_185_747 vdd_d vss_d / DCAP16LVT
XXFILLER_185_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_185_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_186_747 vdd_d vss_d / DCAP16LVT
XXFILLER_186_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_186_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_187_747 vdd_d vss_d / DCAP16LVT
XXFILLER_187_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_187_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_188_747 vdd_d vss_d / DCAP16LVT
XXFILLER_188_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_188_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_189_747 vdd_d vss_d / DCAP16LVT
XXFILLER_189_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_189_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_190_747 vdd_d vss_d / DCAP16LVT
XXFILLER_190_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_190_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_191_747 vdd_d vss_d / DCAP16LVT
XXFILLER_191_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_191_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_192_747 vdd_d vss_d / DCAP16LVT
XXFILLER_192_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_192_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_193_747 vdd_d vss_d / DCAP16LVT
XXFILLER_193_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_193_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_194_747 vdd_d vss_d / DCAP16LVT
XXFILLER_194_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_194_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_195_747 vdd_d vss_d / DCAP16LVT
XXFILLER_195_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_195_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_196_747 vdd_d vss_d / DCAP16LVT
XXFILLER_196_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_196_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_197_747 vdd_d vss_d / DCAP16LVT
XXFILLER_197_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_197_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_198_747 vdd_d vss_d / DCAP16LVT
XXFILLER_198_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_198_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_199_747 vdd_d vss_d / DCAP16LVT
XXFILLER_199_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_199_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_200_747 vdd_d vss_d / DCAP16LVT
XXFILLER_200_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_200_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_201_747 vdd_d vss_d / DCAP16LVT
XXFILLER_201_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_201_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_202_747 vdd_d vss_d / DCAP16LVT
XXFILLER_202_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_202_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_203_747 vdd_d vss_d / DCAP16LVT
XXFILLER_203_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_203_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_204_747 vdd_d vss_d / DCAP16LVT
XXFILLER_204_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_204_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_205_747 vdd_d vss_d / DCAP16LVT
XXFILLER_205_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_205_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_206_416 vdd_d vss_d / DCAP16LVT
XXFILLER_206_927 vdd_d vss_d / DCAP16LVT
XXFILLER_206_1404 vdd_d vss_d / DCAP16LVT
XXFILLER_207_2326 vdd_d vss_d / DCAP16LVT
XXFILLER_214_672 vdd_d vss_d / DCAP16LVT
XXFILLER_214_2321 vdd_d vss_d / DCAP16LVT
XXFILLER_219_2320 vdd_d vss_d / DCAP16LVT
XXFILLER_223_747 vdd_d vss_d / DCAP16LVT
XXFILLER_223_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_223_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_224_747 vdd_d vss_d / DCAP16LVT
XXFILLER_224_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_224_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_225_747 vdd_d vss_d / DCAP16LVT
XXFILLER_225_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_225_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_226_747 vdd_d vss_d / DCAP16LVT
XXFILLER_226_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_226_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_227_747 vdd_d vss_d / DCAP16LVT
XXFILLER_227_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_227_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_228_747 vdd_d vss_d / DCAP16LVT
XXFILLER_228_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_228_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_229_747 vdd_d vss_d / DCAP16LVT
XXFILLER_229_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_229_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_230_747 vdd_d vss_d / DCAP16LVT
XXFILLER_230_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_230_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_231_747 vdd_d vss_d / DCAP16LVT
XXFILLER_231_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_231_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_232_747 vdd_d vss_d / DCAP16LVT
XXFILLER_232_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_232_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_233_747 vdd_d vss_d / DCAP16LVT
XXFILLER_233_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_233_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_234_747 vdd_d vss_d / DCAP16LVT
XXFILLER_234_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_234_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_235_747 vdd_d vss_d / DCAP16LVT
XXFILLER_235_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_235_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_236_747 vdd_d vss_d / DCAP16LVT
XXFILLER_236_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_236_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_237_747 vdd_d vss_d / DCAP16LVT
XXFILLER_237_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_237_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_238_747 vdd_d vss_d / DCAP16LVT
XXFILLER_238_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_238_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_239_747 vdd_d vss_d / DCAP16LVT
XXFILLER_239_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_239_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_240_747 vdd_d vss_d / DCAP16LVT
XXFILLER_240_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_240_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_241_747 vdd_d vss_d / DCAP16LVT
XXFILLER_241_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_241_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_242_747 vdd_d vss_d / DCAP16LVT
XXFILLER_242_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_242_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_243_747 vdd_d vss_d / DCAP16LVT
XXFILLER_243_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_243_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_244_747 vdd_d vss_d / DCAP16LVT
XXFILLER_244_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_244_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_245_747 vdd_d vss_d / DCAP16LVT
XXFILLER_245_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_245_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_246_747 vdd_d vss_d / DCAP16LVT
XXFILLER_246_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_246_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_247_747 vdd_d vss_d / DCAP16LVT
XXFILLER_247_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_247_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_248_747 vdd_d vss_d / DCAP16LVT
XXFILLER_248_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_248_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_249_747 vdd_d vss_d / DCAP16LVT
XXFILLER_249_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_249_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_250_747 vdd_d vss_d / DCAP16LVT
XXFILLER_250_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_250_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_251_747 vdd_d vss_d / DCAP16LVT
XXFILLER_251_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_251_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_252_747 vdd_d vss_d / DCAP16LVT
XXFILLER_252_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_252_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_253_747 vdd_d vss_d / DCAP16LVT
XXFILLER_253_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_253_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_254_747 vdd_d vss_d / DCAP16LVT
XXFILLER_254_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_254_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_255_747 vdd_d vss_d / DCAP16LVT
XXFILLER_255_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_255_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_256_747 vdd_d vss_d / DCAP16LVT
XXFILLER_256_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_256_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_257_747 vdd_d vss_d / DCAP16LVT
XXFILLER_257_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_257_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_258_747 vdd_d vss_d / DCAP16LVT
XXFILLER_258_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_258_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_259_747 vdd_d vss_d / DCAP16LVT
XXFILLER_259_1247 vdd_d vss_d / DCAP16LVT
XXFILLER_259_1747 vdd_d vss_d / DCAP16LVT
XXFILLER_18_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_15_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_14_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_17_512 vdd_d vss_d / DCAP32LVT
XXFILLER_16_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_13_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_12_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_10_768 vdd_d vss_d / DCAP32LVT
XXFILLER_9_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_8_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_7_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_6_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_5_2299 vdd_d vss_d / DCAP32LVT
XXFILLER_1_2303 vdd_d vss_d / DCAP32LVT
XXFILLER_1_768 vdd_d vss_d / DCAP32LVT
XXFILLER_0_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_20_1103 vdd_d vss_d / DCAP32LVT
XXFILLER_19_1122 vdd_d vss_d / DCAP32LVT
XXFILLER_20_1172 vdd_d vss_d / DCAP32LVT
XXFILLER_20_1572 vdd_d vss_d / DCAP32LVT
XXFILLER_21_1110 vdd_d vss_d / DCAP32LVT
XXFILLER_21_1252 vdd_d vss_d / DCAP32LVT
XXFILLER_21_1549 vdd_d vss_d / DCAP32LVT
XXFILLER_21_2318 vdd_d vss_d / DCAP32LVT
XXFILLER_22_1088 vdd_d vss_d / DCAP32LVT
XXFILLER_22_2295 vdd_d vss_d / DCAP32LVT
XXFILLER_23_384 vdd_d vss_d / DCAP32LVT
XXFILLER_23_1315 vdd_d vss_d / DCAP32LVT
XXFILLER_23_2289 vdd_d vss_d / DCAP32LVT
XXFILLER_24_1035 vdd_d vss_d / DCAP32LVT
XXFILLER_24_1620 vdd_d vss_d / DCAP32LVT
XXFILLER_24_2309 vdd_d vss_d / DCAP32LVT
XXFILLER_25_1077 vdd_d vss_d / DCAP32LVT
XXFILLER_25_1177 vdd_d vss_d / DCAP32LVT
XXFILLER_25_1247 vdd_d vss_d / DCAP32LVT
XXFILLER_25_2314 vdd_d vss_d / DCAP32LVT
XXFILLER_26_1374 vdd_d vss_d / DCAP32LVT
XXFILLER_26_1691 vdd_d vss_d / DCAP32LVT
XXFILLER_26_2317 vdd_d vss_d / DCAP32LVT
XXFILLER_27_976 vdd_d vss_d / DCAP32LVT
XXFILLER_27_2288 vdd_d vss_d / DCAP32LVT
XXFILLER_28_384 vdd_d vss_d / DCAP32LVT
XXFILLER_28_862 vdd_d vss_d / DCAP32LVT
XXFILLER_28_1112 vdd_d vss_d / DCAP32LVT
XXFILLER_29_384 vdd_d vss_d / DCAP32LVT
XXFILLER_29_865 vdd_d vss_d / DCAP32LVT
XXFILLER_29_1791 vdd_d vss_d / DCAP32LVT
XXFILLER_29_2303 vdd_d vss_d / DCAP32LVT
XXFILLER_30_384 vdd_d vss_d / DCAP32LVT
XXFILLER_31_1010 vdd_d vss_d / DCAP32LVT
XXFILLER_31_1432 vdd_d vss_d / DCAP32LVT
XXFILLER_31_1816 vdd_d vss_d / DCAP32LVT
XXFILLER_32_748 vdd_d vss_d / DCAP32LVT
XXFILLER_32_934 vdd_d vss_d / DCAP32LVT
XXFILLER_32_1062 vdd_d vss_d / DCAP32LVT
XXFILLER_32_1805 vdd_d vss_d / DCAP32LVT
XXFILLER_32_2310 vdd_d vss_d / DCAP32LVT
XXFILLER_33_384 vdd_d vss_d / DCAP32LVT
XXFILLER_33_1095 vdd_d vss_d / DCAP32LVT
XXFILLER_33_1152 vdd_d vss_d / DCAP32LVT
XXFILLER_33_1225 vdd_d vss_d / DCAP32LVT
XXFILLER_33_1295 vdd_d vss_d / DCAP32LVT
XXFILLER_33_1751 vdd_d vss_d / DCAP32LVT
XXFILLER_34_1035 vdd_d vss_d / DCAP32LVT
XXFILLER_34_1369 vdd_d vss_d / DCAP32LVT
XXFILLER_35_448 vdd_d vss_d / DCAP32LVT
XXFILLER_35_540 vdd_d vss_d / DCAP32LVT
XXFILLER_35_848 vdd_d vss_d / DCAP32LVT
XXFILLER_35_916 vdd_d vss_d / DCAP32LVT
XXFILLER_35_1058 vdd_d vss_d / DCAP32LVT
XXFILLER_35_1259 vdd_d vss_d / DCAP32LVT
XXFILLER_35_1373 vdd_d vss_d / DCAP32LVT
XXFILLER_35_2299 vdd_d vss_d / DCAP32LVT
XXFILLER_36_761 vdd_d vss_d / DCAP32LVT
XXFILLER_36_818 vdd_d vss_d / DCAP32LVT
XXFILLER_36_1530 vdd_d vss_d / DCAP32LVT
XXFILLER_37_493 vdd_d vss_d / DCAP32LVT
XXFILLER_37_738 vdd_d vss_d / DCAP32LVT
XXFILLER_37_1101 vdd_d vss_d / DCAP32LVT
XXFILLER_37_1234 vdd_d vss_d / DCAP32LVT
XXFILLER_37_1417 vdd_d vss_d / DCAP32LVT
XXFILLER_37_1595 vdd_d vss_d / DCAP32LVT
XXFILLER_37_2315 vdd_d vss_d / DCAP32LVT
XXFILLER_38_384 vdd_d vss_d / DCAP32LVT
XXFILLER_38_589 vdd_d vss_d / DCAP32LVT
XXFILLER_38_1395 vdd_d vss_d / DCAP32LVT
XXFILLER_38_1700 vdd_d vss_d / DCAP32LVT
XXFILLER_38_1748 vdd_d vss_d / DCAP32LVT
XXFILLER_38_1886 vdd_d vss_d / DCAP32LVT
XXFILLER_38_2290 vdd_d vss_d / DCAP32LVT
XXFILLER_39_712 vdd_d vss_d / DCAP32LVT
XXFILLER_39_1203 vdd_d vss_d / DCAP32LVT
XXFILLER_39_1784 vdd_d vss_d / DCAP32LVT
XXFILLER_39_2296 vdd_d vss_d / DCAP32LVT
XXFILLER_40_736 vdd_d vss_d / DCAP32LVT
XXFILLER_40_1235 vdd_d vss_d / DCAP32LVT
XXFILLER_40_1307 vdd_d vss_d / DCAP32LVT
XXFILLER_40_1464 vdd_d vss_d / DCAP32LVT
XXFILLER_40_1533 vdd_d vss_d / DCAP32LVT
XXFILLER_40_2317 vdd_d vss_d / DCAP32LVT
XXFILLER_41_768 vdd_d vss_d / DCAP32LVT
XXFILLER_41_890 vdd_d vss_d / DCAP32LVT
XXFILLER_41_1538 vdd_d vss_d / DCAP32LVT
XXFILLER_41_2307 vdd_d vss_d / DCAP32LVT
XXFILLER_42_1287 vdd_d vss_d / DCAP32LVT
XXFILLER_42_1430 vdd_d vss_d / DCAP32LVT
XXFILLER_42_1765 vdd_d vss_d / DCAP32LVT
XXFILLER_42_2296 vdd_d vss_d / DCAP32LVT
XXFILLER_43_1325 vdd_d vss_d / DCAP32LVT
XXFILLER_43_1407 vdd_d vss_d / DCAP32LVT
XXFILLER_43_1562 vdd_d vss_d / DCAP32LVT
XXFILLER_43_1607 vdd_d vss_d / DCAP32LVT
XXFILLER_43_1745 vdd_d vss_d / DCAP32LVT
XXFILLER_43_2306 vdd_d vss_d / DCAP32LVT
XXFILLER_44_320 vdd_d vss_d / DCAP32LVT
XXFILLER_44_842 vdd_d vss_d / DCAP32LVT
XXFILLER_44_954 vdd_d vss_d / DCAP32LVT
XXFILLER_44_1035 vdd_d vss_d / DCAP32LVT
XXFILLER_44_1235 vdd_d vss_d / DCAP32LVT
XXFILLER_44_1313 vdd_d vss_d / DCAP32LVT
XXFILLER_44_1429 vdd_d vss_d / DCAP32LVT
XXFILLER_44_1684 vdd_d vss_d / DCAP32LVT
XXFILLER_45_800 vdd_d vss_d / DCAP32LVT
XXFILLER_45_1528 vdd_d vss_d / DCAP32LVT
XXFILLER_45_1607 vdd_d vss_d / DCAP32LVT
XXFILLER_45_1846 vdd_d vss_d / DCAP32LVT
XXFILLER_45_2291 vdd_d vss_d / DCAP32LVT
XXFILLER_46_1358 vdd_d vss_d / DCAP32LVT
XXFILLER_46_1905 vdd_d vss_d / DCAP32LVT
XXFILLER_46_2303 vdd_d vss_d / DCAP32LVT
XXFILLER_48_882 vdd_d vss_d / DCAP32LVT
XXFILLER_48_2205 vdd_d vss_d / DCAP32LVT
XXFILLER_49_1447 vdd_d vss_d / DCAP32LVT
XXFILLER_49_2289 vdd_d vss_d / DCAP32LVT
XXFILLER_50_763 vdd_d vss_d / DCAP32LVT
XXFILLER_51_1216 vdd_d vss_d / DCAP32LVT
XXFILLER_51_2317 vdd_d vss_d / DCAP32LVT
XXFILLER_52_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_53_1152 vdd_d vss_d / DCAP32LVT
XXFILLER_54_768 vdd_d vss_d / DCAP32LVT
XXFILLER_54_861 vdd_d vss_d / DCAP32LVT
XXFILLER_54_1895 vdd_d vss_d / DCAP32LVT
XXFILLER_55_384 vdd_d vss_d / DCAP32LVT
XXFILLER_55_1904 vdd_d vss_d / DCAP32LVT
XXFILLER_55_2298 vdd_d vss_d / DCAP32LVT
XXFILLER_56_715 vdd_d vss_d / DCAP32LVT
XXFILLER_56_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_56_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_57_715 vdd_d vss_d / DCAP32LVT
XXFILLER_57_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_57_1705 vdd_d vss_d / DCAP32LVT
XXFILLER_58_715 vdd_d vss_d / DCAP32LVT
XXFILLER_58_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_58_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_59_715 vdd_d vss_d / DCAP32LVT
XXFILLER_59_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_59_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_60_715 vdd_d vss_d / DCAP32LVT
XXFILLER_60_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_60_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_61_715 vdd_d vss_d / DCAP32LVT
XXFILLER_61_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_61_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_62_715 vdd_d vss_d / DCAP32LVT
XXFILLER_62_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_62_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_63_715 vdd_d vss_d / DCAP32LVT
XXFILLER_63_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_63_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_64_715 vdd_d vss_d / DCAP32LVT
XXFILLER_64_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_64_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_65_715 vdd_d vss_d / DCAP32LVT
XXFILLER_65_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_65_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_66_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_66_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_67_715 vdd_d vss_d / DCAP32LVT
XXFILLER_67_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_67_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_68_715 vdd_d vss_d / DCAP32LVT
XXFILLER_68_1221 vdd_d vss_d / DCAP32LVT
XXFILLER_68_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_69_192 vdd_d vss_d / DCAP32LVT
XXFILLER_69_715 vdd_d vss_d / DCAP32LVT
XXFILLER_69_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_69_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_69_2295 vdd_d vss_d / DCAP32LVT
XXFILLER_70_715 vdd_d vss_d / DCAP32LVT
XXFILLER_70_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_70_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_71_715 vdd_d vss_d / DCAP32LVT
XXFILLER_71_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_71_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_72_715 vdd_d vss_d / DCAP32LVT
XXFILLER_72_1216 vdd_d vss_d / DCAP32LVT
XXFILLER_72_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_73_192 vdd_d vss_d / DCAP32LVT
XXFILLER_73_715 vdd_d vss_d / DCAP32LVT
XXFILLER_73_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_73_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_73_2314 vdd_d vss_d / DCAP32LVT
XXFILLER_74_715 vdd_d vss_d / DCAP32LVT
XXFILLER_74_1087 vdd_d vss_d / DCAP32LVT
XXFILLER_74_1201 vdd_d vss_d / DCAP32LVT
XXFILLER_74_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_75_715 vdd_d vss_d / DCAP32LVT
XXFILLER_75_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_75_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_76_192 vdd_d vss_d / DCAP32LVT
XXFILLER_76_715 vdd_d vss_d / DCAP32LVT
XXFILLER_76_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_76_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_77_715 vdd_d vss_d / DCAP32LVT
XXFILLER_77_1151 vdd_d vss_d / DCAP32LVT
XXFILLER_77_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_78_715 vdd_d vss_d / DCAP32LVT
XXFILLER_78_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_78_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_79_715 vdd_d vss_d / DCAP32LVT
XXFILLER_79_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_79_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_80_715 vdd_d vss_d / DCAP32LVT
XXFILLER_80_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_80_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_81_715 vdd_d vss_d / DCAP32LVT
XXFILLER_81_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_81_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_82_715 vdd_d vss_d / DCAP32LVT
XXFILLER_82_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_82_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_82_2288 vdd_d vss_d / DCAP32LVT
XXFILLER_83_192 vdd_d vss_d / DCAP32LVT
XXFILLER_83_715 vdd_d vss_d / DCAP32LVT
XXFILLER_83_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_84_715 vdd_d vss_d / DCAP32LVT
XXFILLER_84_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_84_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_85_715 vdd_d vss_d / DCAP32LVT
XXFILLER_85_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_85_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_85_2288 vdd_d vss_d / DCAP32LVT
XXFILLER_86_715 vdd_d vss_d / DCAP32LVT
XXFILLER_86_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_86_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_87_715 vdd_d vss_d / DCAP32LVT
XXFILLER_87_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_87_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_88_715 vdd_d vss_d / DCAP32LVT
XXFILLER_88_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_88_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_89_715 vdd_d vss_d / DCAP32LVT
XXFILLER_89_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_89_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_90_715 vdd_d vss_d / DCAP32LVT
XXFILLER_90_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_90_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_91_715 vdd_d vss_d / DCAP32LVT
XXFILLER_91_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_91_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_92_715 vdd_d vss_d / DCAP32LVT
XXFILLER_92_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_93_715 vdd_d vss_d / DCAP32LVT
XXFILLER_93_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_94_587 vdd_d vss_d / DCAP32LVT
XXFILLER_94_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_94_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_95_1372 vdd_d vss_d / DCAP32LVT
XXFILLER_95_1835 vdd_d vss_d / DCAP32LVT
XXFILLER_96_320 vdd_d vss_d / DCAP32LVT
XXFILLER_96_415 vdd_d vss_d / DCAP32LVT
XXFILLER_96_2292 vdd_d vss_d / DCAP32LVT
XXFILLER_97_2294 vdd_d vss_d / DCAP32LVT
XXFILLER_98_384 vdd_d vss_d / DCAP32LVT
XXFILLER_98_1756 vdd_d vss_d / DCAP32LVT
XXFILLER_99_1374 vdd_d vss_d / DCAP32LVT
XXFILLER_99_1874 vdd_d vss_d / DCAP32LVT
XXFILLER_99_2312 vdd_d vss_d / DCAP32LVT
XXFILLER_100_2296 vdd_d vss_d / DCAP32LVT
XXFILLER_101_1917 vdd_d vss_d / DCAP32LVT
XXFILLER_101_2292 vdd_d vss_d / DCAP32LVT
XXFILLER_102_640 vdd_d vss_d / DCAP32LVT
XXFILLER_102_1134 vdd_d vss_d / DCAP32LVT
XXFILLER_102_1262 vdd_d vss_d / DCAP32LVT
XXFILLER_102_2308 vdd_d vss_d / DCAP32LVT
XXFILLER_103_1719 vdd_d vss_d / DCAP32LVT
XXFILLER_103_1852 vdd_d vss_d / DCAP32LVT
XXFILLER_104_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_105_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_106_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_107_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_109_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_110_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_111_1431 vdd_d vss_d / DCAP32LVT
XXFILLER_111_1809 vdd_d vss_d / DCAP32LVT
XXFILLER_112_715 vdd_d vss_d / DCAP32LVT
XXFILLER_112_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_112_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_113_715 vdd_d vss_d / DCAP32LVT
XXFILLER_113_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_113_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_114_715 vdd_d vss_d / DCAP32LVT
XXFILLER_114_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_114_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_115_715 vdd_d vss_d / DCAP32LVT
XXFILLER_115_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_115_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_116_715 vdd_d vss_d / DCAP32LVT
XXFILLER_116_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_116_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_117_715 vdd_d vss_d / DCAP32LVT
XXFILLER_117_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_117_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_118_715 vdd_d vss_d / DCAP32LVT
XXFILLER_118_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_118_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_119_715 vdd_d vss_d / DCAP32LVT
XXFILLER_119_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_119_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_120_715 vdd_d vss_d / DCAP32LVT
XXFILLER_120_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_120_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_121_715 vdd_d vss_d / DCAP32LVT
XXFILLER_121_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_121_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_122_715 vdd_d vss_d / DCAP32LVT
XXFILLER_122_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_122_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_123_715 vdd_d vss_d / DCAP32LVT
XXFILLER_123_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_123_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_124_715 vdd_d vss_d / DCAP32LVT
XXFILLER_124_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_124_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_125_715 vdd_d vss_d / DCAP32LVT
XXFILLER_125_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_125_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_126_715 vdd_d vss_d / DCAP32LVT
XXFILLER_126_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_126_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_127_715 vdd_d vss_d / DCAP32LVT
XXFILLER_127_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_127_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_128_715 vdd_d vss_d / DCAP32LVT
XXFILLER_128_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_128_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_129_715 vdd_d vss_d / DCAP32LVT
XXFILLER_129_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_129_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_130_715 vdd_d vss_d / DCAP32LVT
XXFILLER_130_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_130_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_131_192 vdd_d vss_d / DCAP32LVT
XXFILLER_131_715 vdd_d vss_d / DCAP32LVT
XXFILLER_131_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_131_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_131_2291 vdd_d vss_d / DCAP32LVT
XXFILLER_132_715 vdd_d vss_d / DCAP32LVT
XXFILLER_132_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_132_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_133_715 vdd_d vss_d / DCAP32LVT
XXFILLER_133_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_133_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_134_715 vdd_d vss_d / DCAP32LVT
XXFILLER_134_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_134_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_135_715 vdd_d vss_d / DCAP32LVT
XXFILLER_135_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_135_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_136_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_136_1587 vdd_d vss_d / DCAP32LVT
XXFILLER_136_1701 vdd_d vss_d / DCAP32LVT
XXFILLER_137_715 vdd_d vss_d / DCAP32LVT
XXFILLER_137_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_137_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_138_715 vdd_d vss_d / DCAP32LVT
XXFILLER_138_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_138_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_139_715 vdd_d vss_d / DCAP32LVT
XXFILLER_139_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_139_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_140_715 vdd_d vss_d / DCAP32LVT
XXFILLER_140_1208 vdd_d vss_d / DCAP32LVT
XXFILLER_140_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_141_715 vdd_d vss_d / DCAP32LVT
XXFILLER_141_1214 vdd_d vss_d / DCAP32LVT
XXFILLER_141_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_142_715 vdd_d vss_d / DCAP32LVT
XXFILLER_142_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_143_715 vdd_d vss_d / DCAP32LVT
XXFILLER_143_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_143_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_144_715 vdd_d vss_d / DCAP32LVT
XXFILLER_144_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_144_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_145_715 vdd_d vss_d / DCAP32LVT
XXFILLER_145_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_145_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_146_715 vdd_d vss_d / DCAP32LVT
XXFILLER_146_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_146_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_147_715 vdd_d vss_d / DCAP32LVT
XXFILLER_147_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_147_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_148_715 vdd_d vss_d / DCAP32LVT
XXFILLER_148_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_148_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_149_715 vdd_d vss_d / DCAP32LVT
XXFILLER_149_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_149_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_150_384 vdd_d vss_d / DCAP32LVT
XXFILLER_150_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_151_384 vdd_d vss_d / DCAP32LVT
XXFILLER_151_904 vdd_d vss_d / DCAP32LVT
XXFILLER_151_1359 vdd_d vss_d / DCAP32LVT
XXFILLER_151_1891 vdd_d vss_d / DCAP32LVT
XXFILLER_151_2318 vdd_d vss_d / DCAP32LVT
XXFILLER_152_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_153_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_154_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_155_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_156_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_157_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_158_640 vdd_d vss_d / DCAP32LVT
XXFILLER_158_2306 vdd_d vss_d / DCAP32LVT
XXFILLER_159_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_160_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_161_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_162_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_163_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_164_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_166_1827 vdd_d vss_d / DCAP32LVT
XXFILLER_167_715 vdd_d vss_d / DCAP32LVT
XXFILLER_167_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_167_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_168_715 vdd_d vss_d / DCAP32LVT
XXFILLER_168_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_168_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_169_715 vdd_d vss_d / DCAP32LVT
XXFILLER_169_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_169_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_170_715 vdd_d vss_d / DCAP32LVT
XXFILLER_170_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_170_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_171_715 vdd_d vss_d / DCAP32LVT
XXFILLER_171_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_171_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_172_715 vdd_d vss_d / DCAP32LVT
XXFILLER_172_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_172_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_173_715 vdd_d vss_d / DCAP32LVT
XXFILLER_173_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_173_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_174_715 vdd_d vss_d / DCAP32LVT
XXFILLER_174_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_174_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_175_715 vdd_d vss_d / DCAP32LVT
XXFILLER_175_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_175_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_176_715 vdd_d vss_d / DCAP32LVT
XXFILLER_176_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_176_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_177_715 vdd_d vss_d / DCAP32LVT
XXFILLER_177_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_177_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_178_715 vdd_d vss_d / DCAP32LVT
XXFILLER_178_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_178_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_179_715 vdd_d vss_d / DCAP32LVT
XXFILLER_179_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_179_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_180_715 vdd_d vss_d / DCAP32LVT
XXFILLER_180_1208 vdd_d vss_d / DCAP32LVT
XXFILLER_180_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_181_715 vdd_d vss_d / DCAP32LVT
XXFILLER_181_1096 vdd_d vss_d / DCAP32LVT
XXFILLER_181_1213 vdd_d vss_d / DCAP32LVT
XXFILLER_181_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_182_715 vdd_d vss_d / DCAP32LVT
XXFILLER_182_1198 vdd_d vss_d / DCAP32LVT
XXFILLER_182_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_183_715 vdd_d vss_d / DCAP32LVT
XXFILLER_183_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_184_715 vdd_d vss_d / DCAP32LVT
XXFILLER_184_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_184_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_185_715 vdd_d vss_d / DCAP32LVT
XXFILLER_185_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_185_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_186_715 vdd_d vss_d / DCAP32LVT
XXFILLER_186_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_186_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_187_715 vdd_d vss_d / DCAP32LVT
XXFILLER_187_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_187_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_188_715 vdd_d vss_d / DCAP32LVT
XXFILLER_188_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_188_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_189_715 vdd_d vss_d / DCAP32LVT
XXFILLER_189_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_189_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_190_715 vdd_d vss_d / DCAP32LVT
XXFILLER_190_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_190_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_191_715 vdd_d vss_d / DCAP32LVT
XXFILLER_191_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_191_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_192_715 vdd_d vss_d / DCAP32LVT
XXFILLER_192_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_192_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_193_715 vdd_d vss_d / DCAP32LVT
XXFILLER_193_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_193_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_194_715 vdd_d vss_d / DCAP32LVT
XXFILLER_194_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_194_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_195_715 vdd_d vss_d / DCAP32LVT
XXFILLER_195_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_195_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_196_715 vdd_d vss_d / DCAP32LVT
XXFILLER_196_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_196_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_197_715 vdd_d vss_d / DCAP32LVT
XXFILLER_197_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_197_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_198_715 vdd_d vss_d / DCAP32LVT
XXFILLER_198_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_198_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_199_715 vdd_d vss_d / DCAP32LVT
XXFILLER_199_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_199_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_200_715 vdd_d vss_d / DCAP32LVT
XXFILLER_200_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_200_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_201_715 vdd_d vss_d / DCAP32LVT
XXFILLER_201_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_201_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_202_715 vdd_d vss_d / DCAP32LVT
XXFILLER_202_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_202_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_203_715 vdd_d vss_d / DCAP32LVT
XXFILLER_203_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_203_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_204_715 vdd_d vss_d / DCAP32LVT
XXFILLER_204_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_204_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_205_715 vdd_d vss_d / DCAP32LVT
XXFILLER_205_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_205_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_206_384 vdd_d vss_d / DCAP32LVT
XXFILLER_206_895 vdd_d vss_d / DCAP32LVT
XXFILLER_207_896 vdd_d vss_d / DCAP32LVT
XXFILLER_207_2294 vdd_d vss_d / DCAP32LVT
XXFILLER_208_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_209_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_210_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_211_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_212_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_213_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_214_640 vdd_d vss_d / DCAP32LVT
XXFILLER_215_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_216_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_217_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_218_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_219_2288 vdd_d vss_d / DCAP32LVT
XXFILLER_220_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_221_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_222_2304 vdd_d vss_d / DCAP32LVT
XXFILLER_223_715 vdd_d vss_d / DCAP32LVT
XXFILLER_223_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_223_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_224_715 vdd_d vss_d / DCAP32LVT
XXFILLER_224_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_224_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_225_715 vdd_d vss_d / DCAP32LVT
XXFILLER_225_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_225_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_226_715 vdd_d vss_d / DCAP32LVT
XXFILLER_226_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_226_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_227_715 vdd_d vss_d / DCAP32LVT
XXFILLER_227_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_227_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_228_715 vdd_d vss_d / DCAP32LVT
XXFILLER_228_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_228_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_229_715 vdd_d vss_d / DCAP32LVT
XXFILLER_229_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_229_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_230_715 vdd_d vss_d / DCAP32LVT
XXFILLER_230_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_230_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_231_715 vdd_d vss_d / DCAP32LVT
XXFILLER_231_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_231_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_232_715 vdd_d vss_d / DCAP32LVT
XXFILLER_232_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_232_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_233_715 vdd_d vss_d / DCAP32LVT
XXFILLER_233_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_233_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_234_715 vdd_d vss_d / DCAP32LVT
XXFILLER_234_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_234_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_235_715 vdd_d vss_d / DCAP32LVT
XXFILLER_235_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_235_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_236_715 vdd_d vss_d / DCAP32LVT
XXFILLER_236_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_236_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_237_715 vdd_d vss_d / DCAP32LVT
XXFILLER_237_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_237_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_238_715 vdd_d vss_d / DCAP32LVT
XXFILLER_238_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_238_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_239_715 vdd_d vss_d / DCAP32LVT
XXFILLER_239_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_239_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_240_715 vdd_d vss_d / DCAP32LVT
XXFILLER_240_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_240_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_241_715 vdd_d vss_d / DCAP32LVT
XXFILLER_241_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_241_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_242_715 vdd_d vss_d / DCAP32LVT
XXFILLER_242_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_242_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_243_715 vdd_d vss_d / DCAP32LVT
XXFILLER_243_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_243_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_244_715 vdd_d vss_d / DCAP32LVT
XXFILLER_244_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_244_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_245_715 vdd_d vss_d / DCAP32LVT
XXFILLER_245_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_245_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_246_715 vdd_d vss_d / DCAP32LVT
XXFILLER_246_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_246_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_247_715 vdd_d vss_d / DCAP32LVT
XXFILLER_247_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_247_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_248_715 vdd_d vss_d / DCAP32LVT
XXFILLER_248_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_248_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_249_715 vdd_d vss_d / DCAP32LVT
XXFILLER_249_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_249_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_250_715 vdd_d vss_d / DCAP32LVT
XXFILLER_250_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_250_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_251_715 vdd_d vss_d / DCAP32LVT
XXFILLER_251_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_251_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_252_715 vdd_d vss_d / DCAP32LVT
XXFILLER_252_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_252_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_253_715 vdd_d vss_d / DCAP32LVT
XXFILLER_253_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_253_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_254_715 vdd_d vss_d / DCAP32LVT
XXFILLER_254_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_254_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_255_715 vdd_d vss_d / DCAP32LVT
XXFILLER_255_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_255_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_256_715 vdd_d vss_d / DCAP32LVT
XXFILLER_256_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_256_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_257_715 vdd_d vss_d / DCAP32LVT
XXFILLER_257_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_257_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_258_715 vdd_d vss_d / DCAP32LVT
XXFILLER_258_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_258_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_259_715 vdd_d vss_d / DCAP32LVT
XXFILLER_259_1215 vdd_d vss_d / DCAP32LVT
XXFILLER_259_1715 vdd_d vss_d / DCAP32LVT
XXFILLER_11_536 vdd_d vss_d / DCAPLVT
XXFILLER_5_2347 vdd_d vss_d / DCAPLVT
XXFILLER_4_392 vdd_d vss_d / DCAPLVT
XXFILLER_4_406 vdd_d vss_d / DCAPLVT
XXFILLER_3_411 vdd_d vss_d / DCAPLVT
XXFILLER_2_534 vdd_d vss_d / DCAPLVT
XXFILLER_1_2347 vdd_d vss_d / DCAPLVT
XXFILLER_1_824 vdd_d vss_d / DCAPLVT
XXFILLER_19_2347 vdd_d vss_d / DCAPLVT
XXFILLER_20_1208 vdd_d vss_d / DCAPLVT
XXFILLER_21_1243 vdd_d vss_d / DCAPLVT
XXFILLER_21_1284 vdd_d vss_d / DCAPLVT
XXFILLER_22_1326 vdd_d vss_d / DCAPLVT
XXFILLER_22_2347 vdd_d vss_d / DCAPLVT
XXFILLER_23_440 vdd_d vss_d / DCAPLVT
XXFILLER_23_1045 vdd_d vss_d / DCAPLVT
XXFILLER_23_1119 vdd_d vss_d / DCAPLVT
XXFILLER_23_1230 vdd_d vss_d / DCAPLVT
XXFILLER_24_1226 vdd_d vss_d / DCAPLVT
XXFILLER_25_1064 vdd_d vss_d / DCAPLVT
XXFILLER_25_1168 vdd_d vss_d / DCAPLVT
XXFILLER_26_396 vdd_d vss_d / DCAPLVT
XXFILLER_26_1047 vdd_d vss_d / DCAPLVT
XXFILLER_26_1073 vdd_d vss_d / DCAPLVT
XXFILLER_27_495 vdd_d vss_d / DCAPLVT
XXFILLER_28_440 vdd_d vss_d / DCAPLVT
XXFILLER_28_512 vdd_d vss_d / DCAPLVT
XXFILLER_28_597 vdd_d vss_d / DCAPLVT
XXFILLER_29_901 vdd_d vss_d / DCAPLVT
XXFILLER_29_1180 vdd_d vss_d / DCAPLVT
XXFILLER_29_2347 vdd_d vss_d / DCAPLVT
XXFILLER_31_384 vdd_d vss_d / DCAPLVT
XXFILLER_31_481 vdd_d vss_d / DCAPLVT
XXFILLER_31_503 vdd_d vss_d / DCAPLVT
XXFILLER_31_1886 vdd_d vss_d / DCAPLVT
XXFILLER_32_414 vdd_d vss_d / DCAPLVT
XXFILLER_32_1423 vdd_d vss_d / DCAPLVT
XXFILLER_32_1473 vdd_d vss_d / DCAPLVT
XXFILLER_32_1511 vdd_d vss_d / DCAPLVT
XXFILLER_32_1853 vdd_d vss_d / DCAPLVT
XXFILLER_33_1143 vdd_d vss_d / DCAPLVT
XXFILLER_33_1257 vdd_d vss_d / DCAPLVT
XXFILLER_33_1415 vdd_d vss_d / DCAPLVT
XXFILLER_33_1457 vdd_d vss_d / DCAPLVT
XXFILLER_33_2347 vdd_d vss_d / DCAPLVT
XXFILLER_34_408 vdd_d vss_d / DCAPLVT
XXFILLER_34_944 vdd_d vss_d / DCAPLVT
XXFILLER_34_1417 vdd_d vss_d / DCAPLVT
XXFILLER_34_1536 vdd_d vss_d / DCAPLVT
XXFILLER_34_2347 vdd_d vss_d / DCAPLVT
XXFILLER_35_484 vdd_d vss_d / DCAPLVT
XXFILLER_35_1550 vdd_d vss_d / DCAPLVT
XXFILLER_35_2347 vdd_d vss_d / DCAPLVT
XXFILLER_36_809 vdd_d vss_d / DCAPLVT
XXFILLER_36_1117 vdd_d vss_d / DCAPLVT
XXFILLER_36_1155 vdd_d vss_d / DCAPLVT
XXFILLER_36_1294 vdd_d vss_d / DCAPLVT
XXFILLER_36_1562 vdd_d vss_d / DCAPLVT
XXFILLER_37_388 vdd_d vss_d / DCAPLVT
XXFILLER_37_537 vdd_d vss_d / DCAPLVT
XXFILLER_37_1149 vdd_d vss_d / DCAPLVT
XXFILLER_37_1203 vdd_d vss_d / DCAPLVT
XXFILLER_37_1373 vdd_d vss_d / DCAPLVT
XXFILLER_37_1683 vdd_d vss_d / DCAPLVT
XXFILLER_37_1916 vdd_d vss_d / DCAPLVT
XXFILLER_37_2347 vdd_d vss_d / DCAPLVT
XXFILLER_38_1029 vdd_d vss_d / DCAPLVT
XXFILLER_38_1237 vdd_d vss_d / DCAPLVT
XXFILLER_38_1357 vdd_d vss_d / DCAPLVT
XXFILLER_38_1812 vdd_d vss_d / DCAPLVT
XXFILLER_39_842 vdd_d vss_d / DCAPLVT
XXFILLER_39_857 vdd_d vss_d / DCAPLVT
XXFILLER_39_1005 vdd_d vss_d / DCAPLVT
XXFILLER_39_1078 vdd_d vss_d / DCAPLVT
XXFILLER_39_1537 vdd_d vss_d / DCAPLVT
XXFILLER_39_1583 vdd_d vss_d / DCAPLVT
XXFILLER_40_437 vdd_d vss_d / DCAPLVT
XXFILLER_40_689 vdd_d vss_d / DCAPLVT
XXFILLER_40_911 vdd_d vss_d / DCAPLVT
XXFILLER_40_942 vdd_d vss_d / DCAPLVT
XXFILLER_40_1058 vdd_d vss_d / DCAPLVT
XXFILLER_40_1169 vdd_d vss_d / DCAPLVT
XXFILLER_40_1771 vdd_d vss_d / DCAPLVT
XXFILLER_40_1854 vdd_d vss_d / DCAPLVT
XXFILLER_41_392 vdd_d vss_d / DCAPLVT
XXFILLER_41_957 vdd_d vss_d / DCAPLVT
XXFILLER_41_1172 vdd_d vss_d / DCAPLVT
XXFILLER_41_1504 vdd_d vss_d / DCAPLVT
XXFILLER_41_2347 vdd_d vss_d / DCAPLVT
XXFILLER_42_566 vdd_d vss_d / DCAPLVT
XXFILLER_42_825 vdd_d vss_d / DCAPLVT
XXFILLER_42_966 vdd_d vss_d / DCAPLVT
XXFILLER_42_1123 vdd_d vss_d / DCAPLVT
XXFILLER_42_1217 vdd_d vss_d / DCAPLVT
XXFILLER_42_1260 vdd_d vss_d / DCAPLVT
XXFILLER_42_1354 vdd_d vss_d / DCAPLVT
XXFILLER_42_2002 vdd_d vss_d / DCAPLVT
XXFILLER_43_1088 vdd_d vss_d / DCAPLVT
XXFILLER_43_1152 vdd_d vss_d / DCAPLVT
XXFILLER_43_1179 vdd_d vss_d / DCAPLVT
XXFILLER_43_1263 vdd_d vss_d / DCAPLVT
XXFILLER_43_1369 vdd_d vss_d / DCAPLVT
XXFILLER_43_1443 vdd_d vss_d / DCAPLVT
XXFILLER_44_485 vdd_d vss_d / DCAPLVT
XXFILLER_44_916 vdd_d vss_d / DCAPLVT
XXFILLER_44_1087 vdd_d vss_d / DCAPLVT
XXFILLER_44_1184 vdd_d vss_d / DCAPLVT
XXFILLER_44_1373 vdd_d vss_d / DCAPLVT
XXFILLER_44_1398 vdd_d vss_d / DCAPLVT
XXFILLER_44_1481 vdd_d vss_d / DCAPLVT
XXFILLER_44_1510 vdd_d vss_d / DCAPLVT
XXFILLER_44_1609 vdd_d vss_d / DCAPLVT
XXFILLER_44_1837 vdd_d vss_d / DCAPLVT
XXFILLER_44_1862 vdd_d vss_d / DCAPLVT
XXFILLER_45_836 vdd_d vss_d / DCAPLVT
XXFILLER_45_1639 vdd_d vss_d / DCAPLVT
XXFILLER_45_2347 vdd_d vss_d / DCAPLVT
XXFILLER_46_1692 vdd_d vss_d / DCAPLVT
XXFILLER_46_2347 vdd_d vss_d / DCAPLVT
XXFILLER_47_668 vdd_d vss_d / DCAPLVT
XXFILLER_48_2347 vdd_d vss_d / DCAPLVT
XXFILLER_50_1489 vdd_d vss_d / DCAPLVT
XXFILLER_50_1918 vdd_d vss_d / DCAPLVT
XXFILLER_53_1200 vdd_d vss_d / DCAPLVT
XXFILLER_54_905 vdd_d vss_d / DCAPLVT
XXFILLER_56_260 vdd_d vss_d / DCAPLVT
XXFILLER_56_2347 vdd_d vss_d / DCAPLVT
XXFILLER_57_260 vdd_d vss_d / DCAPLVT
XXFILLER_57_2347 vdd_d vss_d / DCAPLVT
XXFILLER_58_260 vdd_d vss_d / DCAPLVT
XXFILLER_58_2347 vdd_d vss_d / DCAPLVT
XXFILLER_59_260 vdd_d vss_d / DCAPLVT
XXFILLER_59_2347 vdd_d vss_d / DCAPLVT
XXFILLER_60_260 vdd_d vss_d / DCAPLVT
XXFILLER_60_2347 vdd_d vss_d / DCAPLVT
XXFILLER_61_260 vdd_d vss_d / DCAPLVT
XXFILLER_61_2347 vdd_d vss_d / DCAPLVT
XXFILLER_62_260 vdd_d vss_d / DCAPLVT
XXFILLER_62_2347 vdd_d vss_d / DCAPLVT
XXFILLER_63_260 vdd_d vss_d / DCAPLVT
XXFILLER_63_2347 vdd_d vss_d / DCAPLVT
XXFILLER_64_260 vdd_d vss_d / DCAPLVT
XXFILLER_64_2347 vdd_d vss_d / DCAPLVT
XXFILLER_65_260 vdd_d vss_d / DCAPLVT
XXFILLER_65_2347 vdd_d vss_d / DCAPLVT
XXFILLER_66_260 vdd_d vss_d / DCAPLVT
XXFILLER_66_2347 vdd_d vss_d / DCAPLVT
XXFILLER_67_260 vdd_d vss_d / DCAPLVT
XXFILLER_67_2347 vdd_d vss_d / DCAPLVT
XXFILLER_68_260 vdd_d vss_d / DCAPLVT
XXFILLER_68_2347 vdd_d vss_d / DCAPLVT
XXFILLER_69_244 vdd_d vss_d / DCAPLVT
XXFILLER_69_2347 vdd_d vss_d / DCAPLVT
XXFILLER_70_260 vdd_d vss_d / DCAPLVT
XXFILLER_70_2347 vdd_d vss_d / DCAPLVT
XXFILLER_71_260 vdd_d vss_d / DCAPLVT
XXFILLER_71_2347 vdd_d vss_d / DCAPLVT
XXFILLER_72_260 vdd_d vss_d / DCAPLVT
XXFILLER_72_1260 vdd_d vss_d / DCAPLVT
XXFILLER_72_2347 vdd_d vss_d / DCAPLVT
XXFILLER_74_260 vdd_d vss_d / DCAPLVT
XXFILLER_74_2347 vdd_d vss_d / DCAPLVT
XXFILLER_75_260 vdd_d vss_d / DCAPLVT
XXFILLER_75_2347 vdd_d vss_d / DCAPLVT
XXFILLER_76_2347 vdd_d vss_d / DCAPLVT
XXFILLER_77_260 vdd_d vss_d / DCAPLVT
XXFILLER_77_2347 vdd_d vss_d / DCAPLVT
XXFILLER_78_260 vdd_d vss_d / DCAPLVT
XXFILLER_78_2347 vdd_d vss_d / DCAPLVT
XXFILLER_79_260 vdd_d vss_d / DCAPLVT
XXFILLER_79_2347 vdd_d vss_d / DCAPLVT
XXFILLER_80_260 vdd_d vss_d / DCAPLVT
XXFILLER_80_2347 vdd_d vss_d / DCAPLVT
XXFILLER_81_260 vdd_d vss_d / DCAPLVT
XXFILLER_81_2347 vdd_d vss_d / DCAPLVT
XXFILLER_82_260 vdd_d vss_d / DCAPLVT
XXFILLER_83_2347 vdd_d vss_d / DCAPLVT
XXFILLER_84_260 vdd_d vss_d / DCAPLVT
XXFILLER_84_2347 vdd_d vss_d / DCAPLVT
XXFILLER_85_260 vdd_d vss_d / DCAPLVT
XXFILLER_86_260 vdd_d vss_d / DCAPLVT
XXFILLER_86_2347 vdd_d vss_d / DCAPLVT
XXFILLER_87_260 vdd_d vss_d / DCAPLVT
XXFILLER_87_2347 vdd_d vss_d / DCAPLVT
XXFILLER_88_260 vdd_d vss_d / DCAPLVT
XXFILLER_88_2347 vdd_d vss_d / DCAPLVT
XXFILLER_89_260 vdd_d vss_d / DCAPLVT
XXFILLER_89_2347 vdd_d vss_d / DCAPLVT
XXFILLER_90_260 vdd_d vss_d / DCAPLVT
XXFILLER_90_2347 vdd_d vss_d / DCAPLVT
XXFILLER_91_260 vdd_d vss_d / DCAPLVT
XXFILLER_91_2347 vdd_d vss_d / DCAPLVT
XXFILLER_92_260 vdd_d vss_d / DCAPLVT
XXFILLER_92_2347 vdd_d vss_d / DCAPLVT
XXFILLER_93_260 vdd_d vss_d / DCAPLVT
XXFILLER_93_2347 vdd_d vss_d / DCAPLVT
XXFILLER_94_260 vdd_d vss_d / DCAPLVT
XXFILLER_94_2347 vdd_d vss_d / DCAPLVT
XXFILLER_95_1416 vdd_d vss_d / DCAPLVT
XXFILLER_95_2347 vdd_d vss_d / DCAPLVT
XXFILLER_97_1450 vdd_d vss_d / DCAPLVT
XXFILLER_100_1176 vdd_d vss_d / DCAPLVT
XXFILLER_101_1152 vdd_d vss_d / DCAPLVT
XXFILLER_102_1166 vdd_d vss_d / DCAPLVT
XXFILLER_108_2347 vdd_d vss_d / DCAPLVT
XXFILLER_112_260 vdd_d vss_d / DCAPLVT
XXFILLER_112_2347 vdd_d vss_d / DCAPLVT
XXFILLER_113_260 vdd_d vss_d / DCAPLVT
XXFILLER_113_2347 vdd_d vss_d / DCAPLVT
XXFILLER_114_260 vdd_d vss_d / DCAPLVT
XXFILLER_114_2347 vdd_d vss_d / DCAPLVT
XXFILLER_115_260 vdd_d vss_d / DCAPLVT
XXFILLER_115_2347 vdd_d vss_d / DCAPLVT
XXFILLER_116_260 vdd_d vss_d / DCAPLVT
XXFILLER_116_2347 vdd_d vss_d / DCAPLVT
XXFILLER_117_260 vdd_d vss_d / DCAPLVT
XXFILLER_117_2347 vdd_d vss_d / DCAPLVT
XXFILLER_118_260 vdd_d vss_d / DCAPLVT
XXFILLER_118_2347 vdd_d vss_d / DCAPLVT
XXFILLER_119_260 vdd_d vss_d / DCAPLVT
XXFILLER_119_2347 vdd_d vss_d / DCAPLVT
XXFILLER_120_260 vdd_d vss_d / DCAPLVT
XXFILLER_120_2347 vdd_d vss_d / DCAPLVT
XXFILLER_121_260 vdd_d vss_d / DCAPLVT
XXFILLER_121_2347 vdd_d vss_d / DCAPLVT
XXFILLER_122_260 vdd_d vss_d / DCAPLVT
XXFILLER_122_2347 vdd_d vss_d / DCAPLVT
XXFILLER_123_260 vdd_d vss_d / DCAPLVT
XXFILLER_123_2347 vdd_d vss_d / DCAPLVT
XXFILLER_124_260 vdd_d vss_d / DCAPLVT
XXFILLER_124_2347 vdd_d vss_d / DCAPLVT
XXFILLER_125_260 vdd_d vss_d / DCAPLVT
XXFILLER_125_2347 vdd_d vss_d / DCAPLVT
XXFILLER_126_260 vdd_d vss_d / DCAPLVT
XXFILLER_126_2347 vdd_d vss_d / DCAPLVT
XXFILLER_127_260 vdd_d vss_d / DCAPLVT
XXFILLER_127_2347 vdd_d vss_d / DCAPLVT
XXFILLER_128_260 vdd_d vss_d / DCAPLVT
XXFILLER_128_2347 vdd_d vss_d / DCAPLVT
XXFILLER_129_260 vdd_d vss_d / DCAPLVT
XXFILLER_129_2347 vdd_d vss_d / DCAPLVT
XXFILLER_130_260 vdd_d vss_d / DCAPLVT
XXFILLER_130_2347 vdd_d vss_d / DCAPLVT
XXFILLER_131_248 vdd_d vss_d / DCAPLVT
XXFILLER_131_2347 vdd_d vss_d / DCAPLVT
XXFILLER_132_260 vdd_d vss_d / DCAPLVT
XXFILLER_132_2347 vdd_d vss_d / DCAPLVT
XXFILLER_133_260 vdd_d vss_d / DCAPLVT
XXFILLER_133_2347 vdd_d vss_d / DCAPLVT
XXFILLER_134_260 vdd_d vss_d / DCAPLVT
XXFILLER_134_2347 vdd_d vss_d / DCAPLVT
XXFILLER_135_260 vdd_d vss_d / DCAPLVT
XXFILLER_135_2347 vdd_d vss_d / DCAPLVT
XXFILLER_136_260 vdd_d vss_d / DCAPLVT
XXFILLER_136_760 vdd_d vss_d / DCAPLVT
XXFILLER_136_2347 vdd_d vss_d / DCAPLVT
XXFILLER_137_260 vdd_d vss_d / DCAPLVT
XXFILLER_137_2347 vdd_d vss_d / DCAPLVT
XXFILLER_138_260 vdd_d vss_d / DCAPLVT
XXFILLER_138_2347 vdd_d vss_d / DCAPLVT
XXFILLER_139_260 vdd_d vss_d / DCAPLVT
XXFILLER_139_2347 vdd_d vss_d / DCAPLVT
XXFILLER_140_260 vdd_d vss_d / DCAPLVT
XXFILLER_140_1260 vdd_d vss_d / DCAPLVT
XXFILLER_140_2347 vdd_d vss_d / DCAPLVT
XXFILLER_141_260 vdd_d vss_d / DCAPLVT
XXFILLER_141_2347 vdd_d vss_d / DCAPLVT
XXFILLER_142_260 vdd_d vss_d / DCAPLVT
XXFILLER_142_1167 vdd_d vss_d / DCAPLVT
XXFILLER_142_2347 vdd_d vss_d / DCAPLVT
XXFILLER_143_260 vdd_d vss_d / DCAPLVT
XXFILLER_143_2347 vdd_d vss_d / DCAPLVT
XXFILLER_144_260 vdd_d vss_d / DCAPLVT
XXFILLER_144_2347 vdd_d vss_d / DCAPLVT
XXFILLER_145_260 vdd_d vss_d / DCAPLVT
XXFILLER_145_2347 vdd_d vss_d / DCAPLVT
XXFILLER_146_260 vdd_d vss_d / DCAPLVT
XXFILLER_146_2347 vdd_d vss_d / DCAPLVT
XXFILLER_147_260 vdd_d vss_d / DCAPLVT
XXFILLER_147_2347 vdd_d vss_d / DCAPLVT
XXFILLER_148_260 vdd_d vss_d / DCAPLVT
XXFILLER_148_2347 vdd_d vss_d / DCAPLVT
XXFILLER_149_260 vdd_d vss_d / DCAPLVT
XXFILLER_149_2347 vdd_d vss_d / DCAPLVT
XXFILLER_150_436 vdd_d vss_d / DCAPLVT
XXFILLER_151_1419 vdd_d vss_d / DCAPLVT
XXFILLER_165_1868 vdd_d vss_d / DCAPLVT
XXFILLER_167_260 vdd_d vss_d / DCAPLVT
XXFILLER_167_2347 vdd_d vss_d / DCAPLVT
XXFILLER_168_260 vdd_d vss_d / DCAPLVT
XXFILLER_168_2347 vdd_d vss_d / DCAPLVT
XXFILLER_169_260 vdd_d vss_d / DCAPLVT
XXFILLER_169_2347 vdd_d vss_d / DCAPLVT
XXFILLER_170_260 vdd_d vss_d / DCAPLVT
XXFILLER_170_2347 vdd_d vss_d / DCAPLVT
XXFILLER_171_260 vdd_d vss_d / DCAPLVT
XXFILLER_171_2347 vdd_d vss_d / DCAPLVT
XXFILLER_172_260 vdd_d vss_d / DCAPLVT
XXFILLER_172_2347 vdd_d vss_d / DCAPLVT
XXFILLER_173_260 vdd_d vss_d / DCAPLVT
XXFILLER_173_2347 vdd_d vss_d / DCAPLVT
XXFILLER_174_260 vdd_d vss_d / DCAPLVT
XXFILLER_174_2347 vdd_d vss_d / DCAPLVT
XXFILLER_175_260 vdd_d vss_d / DCAPLVT
XXFILLER_175_2347 vdd_d vss_d / DCAPLVT
XXFILLER_176_260 vdd_d vss_d / DCAPLVT
XXFILLER_176_2347 vdd_d vss_d / DCAPLVT
XXFILLER_177_260 vdd_d vss_d / DCAPLVT
XXFILLER_177_2347 vdd_d vss_d / DCAPLVT
XXFILLER_178_260 vdd_d vss_d / DCAPLVT
XXFILLER_178_2347 vdd_d vss_d / DCAPLVT
XXFILLER_179_260 vdd_d vss_d / DCAPLVT
XXFILLER_179_2347 vdd_d vss_d / DCAPLVT
XXFILLER_180_260 vdd_d vss_d / DCAPLVT
XXFILLER_180_1260 vdd_d vss_d / DCAPLVT
XXFILLER_180_2347 vdd_d vss_d / DCAPLVT
XXFILLER_181_260 vdd_d vss_d / DCAPLVT
XXFILLER_181_1152 vdd_d vss_d / DCAPLVT
XXFILLER_181_2347 vdd_d vss_d / DCAPLVT
XXFILLER_182_260 vdd_d vss_d / DCAPLVT
XXFILLER_182_1242 vdd_d vss_d / DCAPLVT
XXFILLER_182_2347 vdd_d vss_d / DCAPLVT
XXFILLER_183_260 vdd_d vss_d / DCAPLVT
XXFILLER_183_2347 vdd_d vss_d / DCAPLVT
XXFILLER_184_260 vdd_d vss_d / DCAPLVT
XXFILLER_184_2347 vdd_d vss_d / DCAPLVT
XXFILLER_185_260 vdd_d vss_d / DCAPLVT
XXFILLER_185_2347 vdd_d vss_d / DCAPLVT
XXFILLER_186_260 vdd_d vss_d / DCAPLVT
XXFILLER_186_2347 vdd_d vss_d / DCAPLVT
XXFILLER_187_260 vdd_d vss_d / DCAPLVT
XXFILLER_187_2347 vdd_d vss_d / DCAPLVT
XXFILLER_188_260 vdd_d vss_d / DCAPLVT
XXFILLER_188_2347 vdd_d vss_d / DCAPLVT
XXFILLER_189_260 vdd_d vss_d / DCAPLVT
XXFILLER_189_2347 vdd_d vss_d / DCAPLVT
XXFILLER_190_260 vdd_d vss_d / DCAPLVT
XXFILLER_190_2347 vdd_d vss_d / DCAPLVT
XXFILLER_191_260 vdd_d vss_d / DCAPLVT
XXFILLER_191_2347 vdd_d vss_d / DCAPLVT
XXFILLER_192_260 vdd_d vss_d / DCAPLVT
XXFILLER_192_2347 vdd_d vss_d / DCAPLVT
XXFILLER_193_260 vdd_d vss_d / DCAPLVT
XXFILLER_193_2347 vdd_d vss_d / DCAPLVT
XXFILLER_194_260 vdd_d vss_d / DCAPLVT
XXFILLER_194_2347 vdd_d vss_d / DCAPLVT
XXFILLER_195_260 vdd_d vss_d / DCAPLVT
XXFILLER_195_2347 vdd_d vss_d / DCAPLVT
XXFILLER_196_260 vdd_d vss_d / DCAPLVT
XXFILLER_196_2347 vdd_d vss_d / DCAPLVT
XXFILLER_197_260 vdd_d vss_d / DCAPLVT
XXFILLER_197_2347 vdd_d vss_d / DCAPLVT
XXFILLER_198_260 vdd_d vss_d / DCAPLVT
XXFILLER_198_2347 vdd_d vss_d / DCAPLVT
XXFILLER_199_260 vdd_d vss_d / DCAPLVT
XXFILLER_199_2347 vdd_d vss_d / DCAPLVT
XXFILLER_200_260 vdd_d vss_d / DCAPLVT
XXFILLER_200_2347 vdd_d vss_d / DCAPLVT
XXFILLER_201_260 vdd_d vss_d / DCAPLVT
XXFILLER_201_2347 vdd_d vss_d / DCAPLVT
XXFILLER_202_260 vdd_d vss_d / DCAPLVT
XXFILLER_202_2347 vdd_d vss_d / DCAPLVT
XXFILLER_203_260 vdd_d vss_d / DCAPLVT
XXFILLER_203_2347 vdd_d vss_d / DCAPLVT
XXFILLER_204_260 vdd_d vss_d / DCAPLVT
XXFILLER_204_2347 vdd_d vss_d / DCAPLVT
XXFILLER_205_260 vdd_d vss_d / DCAPLVT
XXFILLER_205_2347 vdd_d vss_d / DCAPLVT
XXFILLER_206_1432 vdd_d vss_d / DCAPLVT
XXFILLER_214_700 vdd_d vss_d / DCAPLVT
XXFILLER_223_260 vdd_d vss_d / DCAPLVT
XXFILLER_223_2347 vdd_d vss_d / DCAPLVT
XXFILLER_224_260 vdd_d vss_d / DCAPLVT
XXFILLER_224_2347 vdd_d vss_d / DCAPLVT
XXFILLER_225_260 vdd_d vss_d / DCAPLVT
XXFILLER_225_2347 vdd_d vss_d / DCAPLVT
XXFILLER_226_260 vdd_d vss_d / DCAPLVT
XXFILLER_226_2347 vdd_d vss_d / DCAPLVT
XXFILLER_227_260 vdd_d vss_d / DCAPLVT
XXFILLER_227_2347 vdd_d vss_d / DCAPLVT
XXFILLER_228_260 vdd_d vss_d / DCAPLVT
XXFILLER_228_2347 vdd_d vss_d / DCAPLVT
XXFILLER_229_260 vdd_d vss_d / DCAPLVT
XXFILLER_229_2347 vdd_d vss_d / DCAPLVT
XXFILLER_230_260 vdd_d vss_d / DCAPLVT
XXFILLER_230_2347 vdd_d vss_d / DCAPLVT
XXFILLER_231_260 vdd_d vss_d / DCAPLVT
XXFILLER_231_2347 vdd_d vss_d / DCAPLVT
XXFILLER_232_260 vdd_d vss_d / DCAPLVT
XXFILLER_232_2347 vdd_d vss_d / DCAPLVT
XXFILLER_233_260 vdd_d vss_d / DCAPLVT
XXFILLER_233_2347 vdd_d vss_d / DCAPLVT
XXFILLER_234_260 vdd_d vss_d / DCAPLVT
XXFILLER_234_2347 vdd_d vss_d / DCAPLVT
XXFILLER_235_260 vdd_d vss_d / DCAPLVT
XXFILLER_235_2347 vdd_d vss_d / DCAPLVT
XXFILLER_236_260 vdd_d vss_d / DCAPLVT
XXFILLER_236_2347 vdd_d vss_d / DCAPLVT
XXFILLER_237_260 vdd_d vss_d / DCAPLVT
XXFILLER_237_2347 vdd_d vss_d / DCAPLVT
XXFILLER_238_260 vdd_d vss_d / DCAPLVT
XXFILLER_238_2347 vdd_d vss_d / DCAPLVT
XXFILLER_239_260 vdd_d vss_d / DCAPLVT
XXFILLER_239_2347 vdd_d vss_d / DCAPLVT
XXFILLER_240_260 vdd_d vss_d / DCAPLVT
XXFILLER_240_2347 vdd_d vss_d / DCAPLVT
XXFILLER_241_260 vdd_d vss_d / DCAPLVT
XXFILLER_241_2347 vdd_d vss_d / DCAPLVT
XXFILLER_242_260 vdd_d vss_d / DCAPLVT
XXFILLER_242_2347 vdd_d vss_d / DCAPLVT
XXFILLER_243_260 vdd_d vss_d / DCAPLVT
XXFILLER_243_2347 vdd_d vss_d / DCAPLVT
XXFILLER_244_260 vdd_d vss_d / DCAPLVT
XXFILLER_244_2347 vdd_d vss_d / DCAPLVT
XXFILLER_245_260 vdd_d vss_d / DCAPLVT
XXFILLER_245_2347 vdd_d vss_d / DCAPLVT
XXFILLER_246_260 vdd_d vss_d / DCAPLVT
XXFILLER_246_2347 vdd_d vss_d / DCAPLVT
XXFILLER_247_260 vdd_d vss_d / DCAPLVT
XXFILLER_247_2347 vdd_d vss_d / DCAPLVT
XXFILLER_248_260 vdd_d vss_d / DCAPLVT
XXFILLER_248_2347 vdd_d vss_d / DCAPLVT
XXFILLER_249_260 vdd_d vss_d / DCAPLVT
XXFILLER_249_2347 vdd_d vss_d / DCAPLVT
XXFILLER_250_260 vdd_d vss_d / DCAPLVT
XXFILLER_250_2347 vdd_d vss_d / DCAPLVT
XXFILLER_251_260 vdd_d vss_d / DCAPLVT
XXFILLER_251_2347 vdd_d vss_d / DCAPLVT
XXFILLER_252_260 vdd_d vss_d / DCAPLVT
XXFILLER_252_2347 vdd_d vss_d / DCAPLVT
XXFILLER_253_260 vdd_d vss_d / DCAPLVT
XXFILLER_253_2347 vdd_d vss_d / DCAPLVT
XXFILLER_254_260 vdd_d vss_d / DCAPLVT
XXFILLER_254_2347 vdd_d vss_d / DCAPLVT
XXFILLER_255_260 vdd_d vss_d / DCAPLVT
XXFILLER_255_2347 vdd_d vss_d / DCAPLVT
XXFILLER_256_260 vdd_d vss_d / DCAPLVT
XXFILLER_256_2347 vdd_d vss_d / DCAPLVT
XXFILLER_257_260 vdd_d vss_d / DCAPLVT
XXFILLER_257_2347 vdd_d vss_d / DCAPLVT
XXFILLER_258_260 vdd_d vss_d / DCAPLVT
XXFILLER_258_2347 vdd_d vss_d / DCAPLVT
XXFILLER_259_260 vdd_d vss_d / DCAPLVT
XXFILLER_259_2347 vdd_d vss_d / DCAPLVT
XXwire2891 net2798 vdd_d vss_d net2891 / CKBD3LVT
XXwire2862 net2863 vdd_d vss_d net2862 / CKBD3LVT
XXwire2832 net2833 vdd_d vss_d net2832 / CKBD3LVT
XXwire2856 net2857 vdd_d vss_d net2856 / CKBD3LVT
XXwire2826 net2827 vdd_d vss_d net2826 / CKBD3LVT
XXwire2810 net2811 vdd_d vss_d net2810 / CKBD3LVT
XXwire2771 net2668 vdd_d vss_d net2771 / CKBD3LVT
XXload_slew2769 net2669 vdd_d vss_d net2769 / CKBD3LVT
XXload_slew2768 net2699 vdd_d vss_d net2768 / CKBD3LVT
XXwire2846 net2847 vdd_d vss_d net2846 / CKBD3LVT
XXwire2840 net2841 vdd_d vss_d net2840 / CKBD3LVT
XXwire2816 net2817 vdd_d vss_d net2816 / CKBD3LVT
XXwire2892 net2789 vdd_d vss_d net2892 / BUFFD3LVT
XXwire2893 net2788 vdd_d vss_d net2893 / BUFFD3LVT
XXwire2894 net2787 vdd_d vss_d net2894 / BUFFD3LVT
XXwire2896 adc_comparator_out[15] vdd_d vss_d net2896 / BUFFD3LVT
XXwire2864 net2866 vdd_d vss_d net2864 / BUFFD3LVT
XXload_slew2889 net2661 vdd_d vss_d net2889 / BUFFD3LVT
XXwire2843 net2844 vdd_d vss_d net2843 / BUFFD3LVT
XXwire2859 net2860 vdd_d vss_d net2859 / BUFFD3LVT
XXwire2829 net2830 vdd_d vss_d net2829 / BUFFD3LVT
XXwire2890 net2785 vdd_d vss_d net2890 / BUFFD3LVT
XXwire2888 net2793 vdd_d vss_d net2888 / BUFFD3LVT
XXwire2834 net2836 vdd_d vss_d net2834 / BUFFD3LVT
XXwire2778 spi_bits[155] vdd_d vss_d net2778 / BUFFD3LVT
XXwire2886 net2799 vdd_d vss_d net2886 / BUFFD3LVT
XXwire2887 net2796 vdd_d vss_d net2887 / BUFFD3LVT
XXwire2881 net2579 vdd_d vss_d net2881 / BUFFD3LVT
XXwire2848 net2850 vdd_d vss_d net2848 / BUFFD3LVT
XXwire2818 net2820 vdd_d vss_d net2818 / BUFFD3LVT
XXwire2813 net2814 vdd_d vss_d net2813 / BUFFD3LVT
XXwire2766 net2701 vdd_d vss_d net2766 / BUFFD3LVT
XXwire2895 adc_comparator_out[4] vdd_d vss_d net2895 / CKBD4LVT
XXwire2863 clknet_1_1_leaf_seq_logic vdd_d vss_d net2863 / CKBD4LVT
XXwire2865 net2866 vdd_d vss_d net2865 / CKBD4LVT
XXwire2866 clknet_1_1_leaf_seq_logic vdd_d vss_d net2866 / CKBD4LVT
XXwire2833 clknet_1_1_leaf_seq_samp vdd_d vss_d net2833 / CKBD4LVT
XXwire2842 net2844 vdd_d vss_d net2842 / CKBD4LVT
XXwire2861 net2862 vdd_d vss_d net2861 / CKBD4LVT
XXwire2855 net2856 vdd_d vss_d net2855 / CKBD4LVT
XXwire2857 clknet_1_0_leaf_seq_logic vdd_d vss_d net2857 / CKBD4LVT
XXwire2858 net2860 vdd_d vss_d net2858 / CKBD4LVT
XXwire2860 clknet_1_0_leaf_seq_logic vdd_d vss_d net2860 / CKBD4LVT
XXwire2828 net2830 vdd_d vss_d net2828 / CKBD4LVT
XXwire2825 net2826 vdd_d vss_d net2825 / CKBD4LVT
XXwire2827 clknet_1_0_leaf_seq_samp vdd_d vss_d net2827 / CKBD4LVT
XXwire2831 net2832 vdd_d vss_d net2831 / CKBD4LVT
XXwire2830 clknet_1_0_leaf_seq_samp vdd_d vss_d net2830 / CKBD4LVT
XXwire2870 clknet_0_spi_sclk vdd_d vss_d net2870 / CKBD4LVT
XXwire2874 net2770 vdd_d vss_d net2874 / CKBD4LVT
XXwire2869 net2871 vdd_d vss_d net2869 / CKBD4LVT
XXwire2844 clknet_1_0_leaf_seq_comp vdd_d vss_d net2844 / CKBD4LVT
XXwire2835 net2836 vdd_d vss_d net2835 / CKBD4LVT
XXwire2811 clknet_1_0_leaf_seq_init vdd_d vss_d net2811 / CKBD4LVT
XXwire2814 clknet_1_0_leaf_seq_init vdd_d vss_d net2814 / CKBD4LVT
XXwire2812 net2814 vdd_d vss_d net2812 / CKBD4LVT
XXwire2809 net2810 vdd_d vss_d net2809 / CKBD4LVT
XXwire2770 net2771 vdd_d vss_d net2770 / CKBD4LVT
XXwire2803 adc_comparator_out[11] vdd_d vss_d net2803 / CKBD4LVT
XXwire2805 adc_comparator_out[10] vdd_d vss_d net2805 / CKBD4LVT
XXwire2789 adc_comparator_out[5] vdd_d vss_d net2789 / CKBD4LVT
XXwire2788 adc_comparator_out[6] vdd_d vss_d net2788 / CKBD4LVT
XXwire2787 adc_comparator_out[7] vdd_d vss_d net2787 / CKBD4LVT
XXwire2786 adc_comparator_out[8] vdd_d vss_d net2786 / CKBD4LVT
XXload_slew2780 net2878 vdd_d vss_d net2780 / CKBD4LVT
XXwire2779 net2780 vdd_d vss_d net2779 / CKBD4LVT
XXwire2784 adc_comparator_out[9] vdd_d vss_d net2784 / CKBD4LVT
XXwire2801 adc_comparator_out[12] vdd_d vss_d net2801 / CKBD4LVT
XXwire2767 net2768 vdd_d vss_d net2767 / CKBD4LVT
XXwire2798 adc_comparator_out[13] vdd_d vss_d net2798 / CKBD4LVT
XXload_slew2882 spi_bits[161] vdd_d vss_d net2882 / CKBD4LVT
XXmax_length2871 clknet_0_spi_sclk vdd_d vss_d net2871 / CKBD4LVT
XXwire2849 net2850 vdd_d vss_d net2849 / CKBD4LVT
XXwire2850 clknet_1_1_leaf_seq_comp vdd_d vss_d net2850 / CKBD4LVT
XXwire2847 clknet_1_1_leaf_seq_comp vdd_d vss_d net2847 / CKBD4LVT
XXwire2845 net2846 vdd_d vss_d net2845 / CKBD4LVT
XXwire2841 clknet_1_0_leaf_seq_comp vdd_d vss_d net2841 / CKBD4LVT
XXwire2839 net2840 vdd_d vss_d net2839 / CKBD4LVT
XXwire2836 clknet_1_1_leaf_seq_samp vdd_d vss_d net2836 / CKBD4LVT
XXwire2820 clknet_1_1_leaf_seq_init vdd_d vss_d net2820 / CKBD4LVT
XXwire2819 net2820 vdd_d vss_d net2819 / CKBD4LVT
XXwire2817 clknet_1_1_leaf_seq_init vdd_d vss_d net2817 / CKBD4LVT
XXwire2815 net2816 vdd_d vss_d net2815 / CKBD4LVT
XXwire2763 net2705 vdd_d vss_d net2763 / CKBD4LVT
XXwire2764 net2673 vdd_d vss_d net2764 / CKBD4LVT
XXwire2867 net2868 vdd_d vss_d net2867 / CKBD8LVT
XXwire2823 net2824 vdd_d vss_d net2823 / CKBD8LVT
XXwire2853 net2854 vdd_d vss_d net2853 / CKBD8LVT
XXwire2868 spi_sclk vdd_d vss_d net2868 / BUFFD4LVT
XXwire2824 seq_samp vdd_d vss_d net2824 / BUFFD4LVT
XXclkload2 clknet_4_5_leaf_spi_sclk vdd_d vss_d _unconnected_181 / BUFFD4LVT
XXclkload1 clknet_4_3_leaf_spi_sclk vdd_d vss_d _unconnected_183 / BUFFD4LVT
XXwire2777 net2778 vdd_d vss_d net2777 / BUFFD4LVT
XXwire2792 net2896 vdd_d vss_d net2792 / BUFFD4LVT
XXwire2772 spi_bits[92] vdd_d vss_d net2772 / BUFFD4LVT
XXwire2795 adc_comparator_out[14] vdd_d vss_d net2795 / BUFFD4LVT
XXwire2875 net2767 vdd_d vss_d net2875 / BUFFD4LVT
XXwire2854 seq_logic vdd_d vss_d net2854 / BUFFD4LVT
XXwire2765 net2766 vdd_d vss_d net2765 / BUFFD4LVT
XXhold2873 spi_bits[26] vdd_d vss_d net2873 / DEL4LVT
XXhold2872 spi_bits[3] vdd_d vss_d net2872 / DEL4LVT
XXload_slew2884 spi_bits[157] vdd_d vss_d net2884 / CKBD1LVT
XXload_slew2774 net2877 vdd_d vss_d net2774 / CKBD1LVT
XXload_slew2773 net2883 vdd_d vss_d net2773 / CKBD1LVT
XXload_slew2781 net2879 vdd_d vss_d net2781 / CKBD1LVT
XXload_slew2782 net2880 vdd_d vss_d net2782 / CKBD1LVT
XXload_slew2885 spi_bits[164] vdd_d vss_d net2885 / CKBD1LVT
XXload_slew2883 spi_bits[158] vdd_d vss_d net2883 / CKBD1LVT
XXload_slew2880 spi_bits[150] vdd_d vss_d net2880 / CKBD1LVT
XXload_slew2879 spi_bits[151] vdd_d vss_d net2879 / CKBD1LVT
XXload_slew2878 spi_bits[154] vdd_d vss_d net2878 / CKBD1LVT
XXload_slew2876 spi_bits[159] vdd_d vss_d net2876 / CKBD1LVT
XXload_slew2877 spi_bits[156] vdd_d vss_d net2877 / CKBD1LVT
XXwire2822 net2823 vdd_d vss_d net2822 / BUFFD8LVT
XXclkload0 clknet_4_0_leaf_spi_sclk vdd_d vss_d _unconnected_182 / BUFFD8LVT
XXwire2807 net2808 vdd_d vss_d net2807 / BUFFD8LVT
XXclkload7 clknet_4_15_leaf_spi_sclk vdd_d vss_d _unconnected_188 / BUFFD8LVT
XXwire2852 net2853 vdd_d vss_d net2852 / BUFFD8LVT
XXwire2837 net2838 vdd_d vss_d net2837 / BUFFD8LVT
XXwire2821 net2822 vdd_d vss_d net2821 / BUFFD12LVT
XXwire2851 net2852 vdd_d vss_d net2851 / BUFFD12LVT
XXclkload6 clknet_4_13_leaf_spi_sclk vdd_d vss_d _unconnected_184 / INVD1LVT
XXclkload3 clknet_4_6_leaf_spi_sclk vdd_d vss_d _unconnected_185 / INVD1LVT
XXwire2808 seq_init vdd_d vss_d net2808 / CKBD6LVT
XXwire2791 net2792 vdd_d vss_d net2791 / CKBD6LVT
XXwire2804 net2805 vdd_d vss_d net2804 / CKBD6LVT
XXwire2776 net2777 vdd_d vss_d net2776 / CKBD6LVT
XXwire2775 net2776 vdd_d vss_d net2775 / CKBD6LVT
XXwire2799 net2800 vdd_d vss_d net2799 / CKBD6LVT
XXwire2793 net2794 vdd_d vss_d net2793 / CKBD6LVT
XXwire2802 net2803 vdd_d vss_d net2802 / CKBD6LVT
XXwire2790 net2791 vdd_d vss_d net2790 / CKBD6LVT
XXwire2800 net2801 vdd_d vss_d net2800 / CKBD6LVT
XXwire2785 net2786 vdd_d vss_d net2785 / CKBD6LVT
XXwire2783 net2784 vdd_d vss_d net2783 / CKBD6LVT
XXwire2797 net2891 vdd_d vss_d net2797 / CKBD6LVT
XXwire2794 net2795 vdd_d vss_d net2794 / CKBD6LVT
XXwire2796 net2797 vdd_d vss_d net2796 / CKBD6LVT
XXwire2838 seq_comp vdd_d vss_d net2838 / CKBD6LVT
XXspi_reg_clk_inv_inv_cell_2806 clknet_4_0_leaf_spi_sclk vdd_d vss_d net2806 / 
+ INVD2LVT
.ENDS

************************************************************************
* Library Name: CoRDIA_ADC_01
* Cell Name:    DECAP_UNIT_SHORT
* View Name:    schematic
************************************************************************

.SUBCKT DECAP_UNIT_SHORT VDD VSS
*.PININFO VDD:B VSS:B
XI0[35] VDD VSS / DCAP32
XI0[34] VDD VSS / DCAP32
XI0[33] VDD VSS / DCAP32
XI0[32] VDD VSS / DCAP32
XI0[31] VDD VSS / DCAP32
XI0[30] VDD VSS / DCAP32
XI0[29] VDD VSS / DCAP32
XI0[28] VDD VSS / DCAP32
XI0[27] VDD VSS / DCAP32
XI0[26] VDD VSS / DCAP32
XI0[25] VDD VSS / DCAP32
XI0[24] VDD VSS / DCAP32
XI0[23] VDD VSS / DCAP32
XI0[22] VDD VSS / DCAP32
XI0[21] VDD VSS / DCAP32
XI0[20] VDD VSS / DCAP32
XI0[19] VDD VSS / DCAP32
XI0[18] VDD VSS / DCAP32
XI0[17] VDD VSS / DCAP32
XI0[16] VDD VSS / DCAP32
XI0[15] VDD VSS / DCAP32
XI0[14] VDD VSS / DCAP32
XI0[13] VDD VSS / DCAP32
XI0[12] VDD VSS / DCAP32
XI0[11] VDD VSS / DCAP32
XI0[10] VDD VSS / DCAP32
XI0[9] VDD VSS / DCAP32
XI0[8] VDD VSS / DCAP32
XI0[7] VDD VSS / DCAP32
XI0[6] VDD VSS / DCAP32
XI0[5] VDD VSS / DCAP32
XI0[4] VDD VSS / DCAP32
XI0[3] VDD VSS / DCAP32
XI0[2] VDD VSS / DCAP32
XI0[1] VDD VSS / DCAP32
XI0[0] VDD VSS / DCAP32
XI1[11] VDD VSS / DCAP16
XI1[10] VDD VSS / DCAP16
XI1[9] VDD VSS / DCAP16
XI1[8] VDD VSS / DCAP16
XI1[7] VDD VSS / DCAP16
XI1[6] VDD VSS / DCAP16
XI1[5] VDD VSS / DCAP16
XI1[4] VDD VSS / DCAP16
XI1[3] VDD VSS / DCAP16
XI1[2] VDD VSS / DCAP16
XI1[1] VDD VSS / DCAP16
XI1[0] VDD VSS / DCAP16
.ENDS

************************************************************************
* Library Name: IOlib
* Cell Name:    VSUB_VSS_CUP_pad
* View Name:    schematic
************************************************************************

.SUBCKT VSUB_VSS_CUP_pad VDD VDDPST VSS VSSPST
*.PININFO VDD:B VDDPST:B VSS:B VSSPST:B
XR0 VSS VSUB_DUMMY rm2 l=2u w=4.38u m=1
.ENDS

************************************************************************
* Library Name: frida
* Cell Name:    frida_top
* View Name:    schematic
************************************************************************

.SUBCKT frida_top clk_comp_n_pad clk_comp_p_pad clk_init_n_pad clk_init_p_pad 
+ clk_logic_n_pad clk_logic_p_pad clk_samp_n_pad clk_samp_p_pad comp_out_n_pad 
+ comp_out_p_pad rst_b_pad spi_cs_b_pad spi_sclk_pad spi_sdi_pad spi_sdo_pad 
+ vdd_a vdd_d vdd_dac vdd_io vin_n_pad vin_p_pad vss_a vss_d vss_dac vss_io
*.PININFO clk_comp_n_pad:B clk_comp_p_pad:B clk_init_n_pad:B clk_init_p_pad:B 
*.PININFO clk_logic_n_pad:B clk_logic_p_pad:B clk_samp_n_pad:B 
*.PININFO clk_samp_p_pad:B comp_out_n_pad:B comp_out_p_pad:B rst_b_pad:B 
*.PININFO spi_cs_b_pad:B spi_sclk_pad:B spi_sdi_pad:B spi_sdo_pad:B vdd_a:B 
*.PININFO vdd_d:B vdd_dac:B vdd_io:B vin_n_pad:B vin_p_pad:B vss_a:B vss_d:B 
*.PININFO vss_dac:B vss_io:B
XI8 net6 net6 net6 net111 net112 comp_out_n_pad comp_out_p_pad net2 vdd_io 
+ vss_d vss_io / LVDS_TX_CUP_pad
XI15 net36 net34 clk_logic_n_pad clk_logic_p_pad net2 vdd_io vss_d vss_io / 
+ LVDS_RX_CUP_pad
XI16 net32 net30 clk_comp_n_pad clk_comp_p_pad net2 vdd_io vss_d vss_io / 
+ LVDS_RX_CUP_pad
XI5 net24 net20 clk_samp_n_pad clk_samp_p_pad net2 vdd_io vss_d vss_io / 
+ LVDS_RX_CUP_pad
XI4 net16 net12 clk_init_n_pad clk_init_p_pad net2 vdd_io vss_d vss_io / 
+ LVDS_RX_CUP_pad
XI6 net83 net19 net83 rst_b_pad net19 net83 net2 vdd_io vss_d vss_io net89 
+ net90 / CMOS_IO_CUP_pad
XI12 net3 net4 net3 spi_sdi_pad net4 net3 net2 vdd_io vss_d vss_io net47 net48 
+ / CMOS_IO_CUP_pad
XI10 net13 net23 net13 spi_cs_b_pad net23 net13 net2 vdd_io vss_d vss_io net9 
+ net108 / CMOS_IO_CUP_pad
XI13 net37 net22 net37 spi_sclk_pad net22 net37 net2 vdd_io vss_d vss_io net45 
+ net46 / CMOS_IO_CUP_pad
XI11 net1 net7 net7 spi_sdo_pad net7 net21 net2 vdd_io vss_d vss_io net5 net60 
+ / CMOS_IO_CUP_pad
XI75 net74 vdd_a vss_d vss_a / POWER_CUP_pad
XI21 net8 vdd_dac vss_d vss_dac / POWER_CUP_pad
XI27 net10 vdd_d vss_d vss_d / POWER_CUP_pad
XI14 net2 vdd_io vss_d vss_io / POWER_CUP_pad
XI24 net76 vin_n vin_n_pad net8 vdd_dac vss_d vss_dac / PASSIVE_CUP_pad
XI23 net69 vin_p vin_p_pad net8 vdd_dac vss_d vss_dac / PASSIVE_CUP_pad
XI70 vdd_io vss_io net83 / TIELLVT
XI67 vdd_io vss_io net13 / TIELLVT
XI64 vdd_io vss_io net21 / TIELLVT
XI61 vdd_io vss_io net3 / TIELLVT
XI58 vdd_io vss_io net37 / TIELLVT
XI53 vdd_io vss_io net16 / TIELLVT
XI52 vdd_io vss_io net24 / TIELLVT
XI51 vdd_io vss_io net32 / TIELLVT
XI50 vdd_io vss_io net36 / TIELLVT
XI73 vdd_io vss_io net111 / TIELLVT
XI87 net74 vdd_a vss_d vss_a / GROUND_CUP_pad
XI22 net8 vdd_dac vss_d vss_dac / GROUND_CUP_pad
XI7 net2 vdd_io vss_d vss_io / GROUND_CUP_pad
XI1 net74 vdd_a vss_d vss_a / GROUND_CUP_pad
XI19 net10 vdd_d vss_d vss_d / GROUND_CUP_pad
XI43 net10 vdd_d vss_d vss_d / GROUND_CUP_pad
XI49[0] vdd_a vss_a / DECAP_UNIT
XI49[1] vdd_a vss_a / DECAP_UNIT
XI49[2] vdd_a vss_a / DECAP_UNIT
XI49[3] vdd_a vss_a / DECAP_UNIT
XI49[4] vdd_a vss_a / DECAP_UNIT
XI49[5] vdd_a vss_a / DECAP_UNIT
XI49[6] vdd_a vss_a / DECAP_UNIT
XI49[7] vdd_a vss_a / DECAP_UNIT
XI49[8] vdd_a vss_a / DECAP_UNIT
XI49[9] vdd_a vss_a / DECAP_UNIT
XI49[10] vdd_a vss_a / DECAP_UNIT
XI49[11] vdd_a vss_a / DECAP_UNIT
XI49[12] vdd_a vss_a / DECAP_UNIT
XI49[13] vdd_a vss_a / DECAP_UNIT
XI49[14] vdd_a vss_a / DECAP_UNIT
XI77[0] vdd_d vss_d / DECAP_UNIT
XI77[1] vdd_d vss_d / DECAP_UNIT
XI77[2] vdd_d vss_d / DECAP_UNIT
XI77[3] vdd_d vss_d / DECAP_UNIT
XI77[4] vdd_d vss_d / DECAP_UNIT
XI77[5] vdd_d vss_d / DECAP_UNIT
XI77[6] vdd_d vss_d / DECAP_UNIT
XI77[7] vdd_d vss_d / DECAP_UNIT
XI77[8] vdd_d vss_d / DECAP_UNIT
XI77[9] vdd_d vss_d / DECAP_UNIT
XI77[10] vdd_d vss_d / DECAP_UNIT
XI77[11] vdd_d vss_d / DECAP_UNIT
XI77[12] vdd_d vss_d / DECAP_UNIT
XI77[13] vdd_d vss_d / DECAP_UNIT
XI77[14] vdd_d vss_d / DECAP_UNIT
XI95 vdd_io vss_io net18 / TIEHLVT
XI94 vdd_io vss_io net17 / TIEHLVT
XI91 vdd_io vss_io net15 / TIEHLVT
XI71 vdd_io vss_io net19 / TIEHLVT
XI66 vdd_io vss_io net23 / TIEHLVT
XI65 vdd_io vss_io net7 / TIEHLVT
XI60 vdd_io vss_io net4 / TIEHLVT
XI57 vdd_io vss_io net22 / TIEHLVT
XI74 vdd_io vss_io net6 / TIEHLVT
XI90 vdd_io vss_io net14 / TIEHLVT
XI98 net112 net89 net30 net12 net34 net20 net9 net45 net47 net1 vdd_a vdd_d 
+ vdd_dac vin_n vin_p vss_a vss_d vss_dac / frida_core
XI78[0] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI78[1] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI78[2] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI78[3] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI78[4] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI78[5] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI78[6] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI78[7] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI78[8] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI78[9] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI78[10] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI78[11] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI78[12] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI78[13] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI78[14] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI78[15] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI78[16] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI78[17] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI78[18] vdd_dac vss_dac / DECAP_UNIT_SHORT
XI79[0] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[1] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[2] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[3] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[4] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[5] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[6] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[7] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[8] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[9] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[10] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[11] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[12] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[13] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[14] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[15] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[16] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[17] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[18] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[19] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[20] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[21] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[22] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[23] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[24] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[25] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[26] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[27] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[28] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[29] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[30] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[31] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[32] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[33] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[34] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[35] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[36] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[37] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[38] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[39] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[40] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[41] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[42] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[43] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[44] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[45] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[46] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[47] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[48] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[49] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[50] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[51] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[52] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[53] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[54] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[55] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[56] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[57] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[58] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[59] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[60] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[61] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[62] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[63] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[64] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[65] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[66] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[67] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[68] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[69] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[70] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[71] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[72] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[73] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[74] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[75] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[76] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[77] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[78] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[79] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[80] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[81] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[82] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[83] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[84] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[85] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[86] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[87] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[88] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[89] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[90] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[91] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[92] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[93] vdd_io vss_io / DECAP_UNIT_SHORT
XI79[94] vdd_io vss_io / DECAP_UNIT_SHORT
XI44 net10 vdd_d vss_d vss_d / VSUB_VSS_CUP_pad
.ENDS

