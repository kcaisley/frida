**********************************************************************

.SUBCKT SARCMPHX1_EV CI CK CO VMR N1 N2 AVDD AVSS
MN0  N1 CK AVSS AVSS NCHDL
MN1  N2 CI N1   AVSS NCHDL
MN2  N1 CI N2   AVSS NCHDL
MN3  N2 CI N1   AVSS NCHDL
MN4  N1 CI N2   AVSS NCHDL
MN5  N2 CI N1   AVSS NCHDL
MN6  CO VMR N2   AVSS NCHDL

MP0  AVDD CK N1 AVDD PCHDL
MP1  N2 CK AVDD AVDD PCHDL
MP2  AVDD AVDD N2 AVDD PCHDL
MP3  CO CK AVDD AVDD PCHDL
MP4  AVDD VMR CO AVDD PCHDL
MP5  CO VMR AVDD AVDD PCHDL
MP6  AVDD VMR CO AVDD PCHDL
.ENDS SARCMPHX1_EV

.SUBCKT SARKICKHX1_EV CI CK CKN AVDD AVSS
MN0  N1 CKN AVSS AVSS NCHDL
MN1  N1 CI N1   AVSS NCHDL
MN2  N1 CI N1   AVSS NCHDL
MN3  N1 CI N1   AVSS NCHDL
MN4  N1 CI N1   AVSS NCHDL
MN5  N1 CI N1   AVSS NCHDL
MN6  AVDD CK N1   AVSS NCHDL

MP0  AVDD CKN N1 AVDD PCHDL
MP1_DMY AVDD AVDD AVDD AVDD PCHDL
MP2_DMY AVDD AVDD AVDD AVDD PCHDL
MP3_DMY AVDD AVDD AVDD AVDD PCHDL
MP4_DMY AVDD AVDD AVDD AVDD PCHDL
MP5_DMY AVDD AVDD AVDD AVDD PCHDL
MP6  AVDD AVDD AVDD AVDD PCHDL
.ENDS SARKICKHX1_EV

.SUBCKT SARCMPX1_EV CPI CNI CPO CNO CK_CMP CK_SAMPLE DONE AVDD AVSS
XA0 AVSS AVDD TAPCELLB_EV
XA1 CPI CK_B CK_N AVDD AVSS SARKICKHX1_EV
XA2 CPI CK_B CNO_I CPO_I N1 NC1 AVDD AVSS SARCMPHX1_EV
XA2a CPO_I CPO AVDD AVSS IVX4_EV
XA3a CNO_I CNO AVDD AVSS IVX4_EV
XA3 CNI CK_B CPO_I CNO_I N1 NC2 AVDD AVSS SARCMPHX1_EV
XA4 CNI CK_B CK_N AVDD AVSS SARKICKHX1_EV
XA9 CK_N CK_B AVDD AVSS IVX1_EV
XA10 DONE_N CK_A CK_N AVDD AVSS NDX1_EV
XA11 CK_SAMPLE DONE DONE_N AVDD AVSS NRX1_EV
XA12 CK_CMP CK_A AVDD AVSS IVX1_EV
XA13 AVSS AVDD TAPCELLB_EV
.ENDS