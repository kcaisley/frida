VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO s
  CLASS COVER ;
  ORIGIN 0 0 ;
  SIZE 5 BY 5 ;
END s

END LIBRARY