* Comparator Topology Netlists
* Figure 4.13(d): Self-timed Double-tail Comparator

* ========================================================================
* (d) Self-timed Double-tail Comparator
* ========================================================================
.SUBCKT comp_selftimed_doubletail in_p in_n out_p out_n clk clk_b vdd_a vss_a
*.PININFO in_p:I in_n:I out_p:O out_n:O clk:I clk_b:I vdd_a:B vss_a:B

* First stage (input stage)
* Tail transistor
MNtail1 tail1 clk vss_a vss_a nmos

* Input differential pair
MNinn xn in_n tail1 vss_a nmos
MNinp xp in_p tail1 vss_a nmos

* First stage intermediate nodes
MNxn midn xn vss_a vss_a nmos
MNxp midp xp vss_a vss_a nmos

* First stage PMOS loads
MPldMN midn xp vdd_a vdd_a pmos
MPldMP midp xn vdd_a vdd_a pmos

* Reset switches for intermediate nodes
MPswMN xn clk vdd_a vdd_a pmos
MPswMP xp clk vdd_a vdd_a pmos

* Second stage
* Tail control (self-timed from first stage)
MNtail2 tail2 midn vss_a vss_a nmos
MNtail2b tail2 midp vss_a vss_a nmos

* Cross-coupled NMOS pair driven by first stage
MNnfbn out_p out_n midp tail2 nmos
MNnfbp out_n out_p midn tail2 nmos

* Output reset switches
MPswon out_n clk vdd_a vdd_a pmos
MPswop out_p clk vdd_a vdd_a pmos

* Cross-coupled PMOS latch
MPpfbn out_n out_p vdd_a vdd_a pmos
MPpfbp out_p out_n vdd_a vdd_a pmos

.ENDS comp_selftimed_doubletail
