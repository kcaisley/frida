// Verilog HDL for "basic", "cds_alias" "functional"

module cds_alias(a,a);
  parameter width = 1;
  inout [width-1:0] a;
endmodule
