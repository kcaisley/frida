module cds_thru(src,dst);
inout src,dst;
    cds_thrualias i0 (src,dst);
endmodule
